
module DELAY_LINE ( RESET, CLK, Delay_Line_in, Delay_Line_address, 
        Delay_Line_sample_shift, Delay_Line_out );
  input [7:0] Delay_Line_in;
  input [4:0] Delay_Line_address;
  output [7:0] Delay_Line_out;
  input RESET, CLK, Delay_Line_sample_shift;
  wire   N2, N3, N4, N5, N6, \x[0][7] , \x[0][6] , \x[0][5] , \x[0][4] ,
         \x[0][3] , \x[0][2] , \x[0][1] , \x[0][0] , \x[1][7] , \x[1][6] ,
         \x[1][5] , \x[1][4] , \x[1][3] , \x[1][2] , \x[1][1] , \x[1][0] ,
         \x[2][7] , \x[2][6] , \x[2][5] , \x[2][4] , \x[2][3] , \x[2][2] ,
         \x[2][1] , \x[2][0] , \x[3][7] , \x[3][6] , \x[3][5] , \x[3][4] ,
         \x[3][3] , \x[3][2] , \x[3][1] , \x[3][0] , \x[4][7] , \x[4][6] ,
         \x[4][5] , \x[4][4] , \x[4][3] , \x[4][2] , \x[4][1] , \x[4][0] ,
         \x[5][7] , \x[5][6] , \x[5][5] , \x[5][4] , \x[5][3] , \x[5][2] ,
         \x[5][1] , \x[5][0] , \x[6][7] , \x[6][6] , \x[6][5] , \x[6][4] ,
         \x[6][3] , \x[6][2] , \x[6][1] , \x[6][0] , \x[7][7] , \x[7][6] ,
         \x[7][5] , \x[7][4] , \x[7][3] , \x[7][2] , \x[7][1] , \x[7][0] ,
         \x[8][7] , \x[8][6] , \x[8][5] , \x[8][4] , \x[8][3] , \x[8][2] ,
         \x[8][1] , \x[8][0] , \x[9][7] , \x[9][6] , \x[9][5] , \x[9][4] ,
         \x[9][3] , \x[9][2] , \x[9][1] , \x[9][0] , \x[10][7] , \x[10][6] ,
         \x[10][5] , \x[10][4] , \x[10][3] , \x[10][2] , \x[10][1] ,
         \x[10][0] , \x[11][7] , \x[11][6] , \x[11][5] , \x[11][4] ,
         \x[11][3] , \x[11][2] , \x[11][1] , \x[11][0] , \x[12][7] ,
         \x[12][6] , \x[12][5] , \x[12][4] , \x[12][3] , \x[12][2] ,
         \x[12][1] , \x[12][0] , \x[13][7] , \x[13][6] , \x[13][5] ,
         \x[13][4] , \x[13][3] , \x[13][2] , \x[13][1] , \x[13][0] ,
         \x[14][7] , \x[14][6] , \x[14][5] , \x[14][4] , \x[14][3] ,
         \x[14][2] , \x[14][1] , \x[14][0] , \x[15][7] , \x[15][6] ,
         \x[15][5] , \x[15][4] , \x[15][3] , \x[15][2] , \x[15][1] ,
         \x[15][0] , \x[16][7] , \x[16][6] , \x[16][5] , \x[16][4] ,
         \x[16][3] , \x[16][2] , \x[16][1] , \x[16][0] , \x[17][7] ,
         \x[17][6] , \x[17][5] , \x[17][4] , \x[17][3] , \x[17][2] ,
         \x[17][1] , \x[17][0] , \x[18][7] , \x[18][6] , \x[18][5] ,
         \x[18][4] , \x[18][3] , \x[18][2] , \x[18][1] , \x[18][0] ,
         \x[19][7] , \x[19][6] , \x[19][5] , \x[19][4] , \x[19][3] ,
         \x[19][2] , \x[19][1] , \x[19][0] , \x[20][7] , \x[20][6] ,
         \x[20][5] , \x[20][4] , \x[20][3] , \x[20][2] , \x[20][1] ,
         \x[20][0] , \x[21][7] , \x[21][6] , \x[21][5] , \x[21][4] ,
         \x[21][3] , \x[21][2] , \x[21][1] , \x[21][0] , \x[22][7] ,
         \x[22][6] , \x[22][5] , \x[22][4] , \x[22][3] , \x[22][2] ,
         \x[22][1] , \x[22][0] , \x[23][7] , \x[23][6] , \x[23][5] ,
         \x[23][4] , \x[23][3] , \x[23][2] , \x[23][1] , \x[23][0] ,
         \x[24][7] , \x[24][6] , \x[24][5] , \x[24][4] , \x[24][3] ,
         \x[24][2] , \x[24][1] , \x[24][0] , \x[25][7] , \x[25][6] ,
         \x[25][5] , \x[25][4] , \x[25][3] , \x[25][2] , \x[25][1] ,
         \x[25][0] , \x[26][7] , \x[26][6] , \x[26][5] , \x[26][4] ,
         \x[26][3] , \x[26][2] , \x[26][1] , \x[26][0] , \x[27][7] ,
         \x[27][6] , \x[27][5] , \x[27][4] , \x[27][3] , \x[27][2] ,
         \x[27][1] , \x[27][0] , \x[28][7] , \x[28][6] , \x[28][5] ,
         \x[28][4] , \x[28][3] , \x[28][2] , \x[28][1] , \x[28][0] ,
         \x[29][7] , \x[29][6] , \x[29][5] , \x[29][4] , \x[29][3] ,
         \x[29][2] , \x[29][1] , \x[29][0] , \x[30][7] , \x[30][6] ,
         \x[30][5] , \x[30][4] , \x[30][3] , \x[30][2] , \x[30][1] ,
         \x[30][0] , \x[31][7] , \x[31][6] , \x[31][5] , \x[31][4] ,
         \x[31][3] , \x[31][2] , \x[31][1] , \x[31][0] , n249, n250, n251,
         n252, n253, n254, n255, n256, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n257, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644;
  assign N2 = Delay_Line_address[0];
  assign N3 = Delay_Line_address[1];
  assign N4 = Delay_Line_address[2];
  assign N5 = Delay_Line_address[3];
  assign N6 = Delay_Line_address[4];

  OAI212 U3 ( .A(n111), .B(n256), .C(n258), .Q(n516) );
  OAI212 U5 ( .A(n112), .B(n255), .C(n260), .Q(n517) );
  OAI212 U7 ( .A(n111), .B(n254), .C(n261), .Q(n518) );
  OAI212 U9 ( .A(n113), .B(n253), .C(n262), .Q(n519) );
  OAI212 U11 ( .A(n113), .B(n252), .C(n263), .Q(n520) );
  OAI212 U13 ( .A(n113), .B(n251), .C(n264), .Q(n521) );
  OAI212 U15 ( .A(n113), .B(n250), .C(n265), .Q(n522) );
  OAI212 U17 ( .A(n113), .B(n249), .C(n266), .Q(n523) );
  DF3 \x_reg[0][7]  ( .D(n644), .C(CLK), .Q(\x[0][7] ) );
  DF3 \x_reg[0][6]  ( .D(n643), .C(CLK), .Q(\x[0][6] ) );
  DF3 \x_reg[0][5]  ( .D(n642), .C(CLK), .Q(\x[0][5] ) );
  DF3 \x_reg[0][4]  ( .D(n641), .C(CLK), .Q(\x[0][4] ) );
  DF3 \x_reg[0][3]  ( .D(n640), .C(CLK), .Q(\x[0][3] ) );
  DF3 \x_reg[0][2]  ( .D(n639), .C(CLK), .Q(\x[0][2] ) );
  DF3 \x_reg[0][1]  ( .D(n638), .C(CLK), .Q(\x[0][1] ) );
  DF3 \x_reg[0][0]  ( .D(n637), .C(CLK), .Q(\x[0][0] ) );
  DF3 \x_reg[1][7]  ( .D(n636), .C(CLK), .Q(\x[1][7] ) );
  DF3 \x_reg[1][6]  ( .D(n635), .C(CLK), .Q(\x[1][6] ) );
  DF3 \x_reg[1][5]  ( .D(n634), .C(CLK), .Q(\x[1][5] ) );
  DF3 \x_reg[1][4]  ( .D(n633), .C(CLK), .Q(\x[1][4] ) );
  DF3 \x_reg[1][3]  ( .D(n632), .C(CLK), .Q(\x[1][3] ) );
  DF3 \x_reg[1][2]  ( .D(n631), .C(CLK), .Q(\x[1][2] ) );
  DF3 \x_reg[1][1]  ( .D(n630), .C(CLK), .Q(\x[1][1] ) );
  DF3 \x_reg[1][0]  ( .D(n629), .C(CLK), .Q(\x[1][0] ) );
  DF3 \x_reg[2][7]  ( .D(n628), .C(CLK), .Q(\x[2][7] ) );
  DF3 \x_reg[2][6]  ( .D(n627), .C(CLK), .Q(\x[2][6] ) );
  DF3 \x_reg[2][5]  ( .D(n626), .C(CLK), .Q(\x[2][5] ) );
  DF3 \x_reg[2][4]  ( .D(n625), .C(CLK), .Q(\x[2][4] ) );
  DF3 \x_reg[2][3]  ( .D(n624), .C(CLK), .Q(\x[2][3] ) );
  DF3 \x_reg[2][2]  ( .D(n623), .C(CLK), .Q(\x[2][2] ) );
  DF3 \x_reg[2][1]  ( .D(n622), .C(CLK), .Q(\x[2][1] ) );
  DF3 \x_reg[2][0]  ( .D(n621), .C(CLK), .Q(\x[2][0] ) );
  DF3 \x_reg[3][7]  ( .D(n620), .C(CLK), .Q(\x[3][7] ) );
  DF3 \x_reg[3][6]  ( .D(n619), .C(CLK), .Q(\x[3][6] ) );
  DF3 \x_reg[3][5]  ( .D(n618), .C(CLK), .Q(\x[3][5] ) );
  DF3 \x_reg[3][4]  ( .D(n617), .C(CLK), .Q(\x[3][4] ) );
  DF3 \x_reg[3][3]  ( .D(n616), .C(CLK), .Q(\x[3][3] ) );
  DF3 \x_reg[3][2]  ( .D(n615), .C(CLK), .Q(\x[3][2] ) );
  DF3 \x_reg[3][1]  ( .D(n614), .C(CLK), .Q(\x[3][1] ) );
  DF3 \x_reg[3][0]  ( .D(n613), .C(CLK), .Q(\x[3][0] ) );
  DF3 \x_reg[4][7]  ( .D(n612), .C(CLK), .Q(\x[4][7] ) );
  DF3 \x_reg[4][6]  ( .D(n611), .C(CLK), .Q(\x[4][6] ) );
  DF3 \x_reg[4][5]  ( .D(n610), .C(CLK), .Q(\x[4][5] ) );
  DF3 \x_reg[4][4]  ( .D(n609), .C(CLK), .Q(\x[4][4] ) );
  DF3 \x_reg[4][3]  ( .D(n608), .C(CLK), .Q(\x[4][3] ) );
  DF3 \x_reg[4][2]  ( .D(n607), .C(CLK), .Q(\x[4][2] ) );
  DF3 \x_reg[4][1]  ( .D(n606), .C(CLK), .Q(\x[4][1] ) );
  DF3 \x_reg[4][0]  ( .D(n605), .C(CLK), .Q(\x[4][0] ) );
  DF3 \x_reg[5][7]  ( .D(n604), .C(CLK), .Q(\x[5][7] ) );
  DF3 \x_reg[5][6]  ( .D(n603), .C(CLK), .Q(\x[5][6] ) );
  DF3 \x_reg[5][5]  ( .D(n602), .C(CLK), .Q(\x[5][5] ) );
  DF3 \x_reg[5][4]  ( .D(n601), .C(CLK), .Q(\x[5][4] ) );
  DF3 \x_reg[5][3]  ( .D(n600), .C(CLK), .Q(\x[5][3] ) );
  DF3 \x_reg[5][2]  ( .D(n599), .C(CLK), .Q(\x[5][2] ) );
  DF3 \x_reg[5][1]  ( .D(n598), .C(CLK), .Q(\x[5][1] ) );
  DF3 \x_reg[5][0]  ( .D(n597), .C(CLK), .Q(\x[5][0] ) );
  DF3 \x_reg[6][7]  ( .D(n596), .C(CLK), .Q(\x[6][7] ) );
  DF3 \x_reg[6][6]  ( .D(n595), .C(CLK), .Q(\x[6][6] ) );
  DF3 \x_reg[6][5]  ( .D(n594), .C(CLK), .Q(\x[6][5] ) );
  DF3 \x_reg[6][4]  ( .D(n593), .C(CLK), .Q(\x[6][4] ) );
  DF3 \x_reg[6][3]  ( .D(n592), .C(CLK), .Q(\x[6][3] ) );
  DF3 \x_reg[6][2]  ( .D(n591), .C(CLK), .Q(\x[6][2] ) );
  DF3 \x_reg[6][1]  ( .D(n590), .C(CLK), .Q(\x[6][1] ) );
  DF3 \x_reg[6][0]  ( .D(n589), .C(CLK), .Q(\x[6][0] ) );
  DF3 \x_reg[7][7]  ( .D(n588), .C(CLK), .Q(\x[7][7] ) );
  DF3 \x_reg[7][6]  ( .D(n587), .C(CLK), .Q(\x[7][6] ) );
  DF3 \x_reg[7][5]  ( .D(n586), .C(CLK), .Q(\x[7][5] ) );
  DF3 \x_reg[7][4]  ( .D(n585), .C(CLK), .Q(\x[7][4] ) );
  DF3 \x_reg[7][3]  ( .D(n584), .C(CLK), .Q(\x[7][3] ) );
  DF3 \x_reg[7][2]  ( .D(n583), .C(CLK), .Q(\x[7][2] ) );
  DF3 \x_reg[7][1]  ( .D(n582), .C(CLK), .Q(\x[7][1] ) );
  DF3 \x_reg[7][0]  ( .D(n581), .C(CLK), .Q(\x[7][0] ) );
  DF3 \x_reg[8][7]  ( .D(n580), .C(CLK), .Q(\x[8][7] ) );
  DF3 \x_reg[8][6]  ( .D(n579), .C(CLK), .Q(\x[8][6] ) );
  DF3 \x_reg[8][5]  ( .D(n578), .C(CLK), .Q(\x[8][5] ) );
  DF3 \x_reg[8][4]  ( .D(n577), .C(CLK), .Q(\x[8][4] ) );
  DF3 \x_reg[8][3]  ( .D(n576), .C(CLK), .Q(\x[8][3] ) );
  DF3 \x_reg[8][2]  ( .D(n575), .C(CLK), .Q(\x[8][2] ) );
  DF3 \x_reg[8][1]  ( .D(n574), .C(CLK), .Q(\x[8][1] ) );
  DF3 \x_reg[8][0]  ( .D(n573), .C(CLK), .Q(\x[8][0] ) );
  DF3 \x_reg[9][7]  ( .D(n572), .C(CLK), .Q(\x[9][7] ) );
  DF3 \x_reg[9][6]  ( .D(n571), .C(CLK), .Q(\x[9][6] ) );
  DF3 \x_reg[9][5]  ( .D(n570), .C(CLK), .Q(\x[9][5] ) );
  DF3 \x_reg[9][4]  ( .D(n569), .C(CLK), .Q(\x[9][4] ) );
  DF3 \x_reg[9][3]  ( .D(n568), .C(CLK), .Q(\x[9][3] ) );
  DF3 \x_reg[9][2]  ( .D(n567), .C(CLK), .Q(\x[9][2] ) );
  DF3 \x_reg[9][1]  ( .D(n566), .C(CLK), .Q(\x[9][1] ) );
  DF3 \x_reg[9][0]  ( .D(n565), .C(CLK), .Q(\x[9][0] ) );
  DF3 \x_reg[10][7]  ( .D(n564), .C(CLK), .Q(\x[10][7] ) );
  DF3 \x_reg[10][6]  ( .D(n563), .C(CLK), .Q(\x[10][6] ) );
  DF3 \x_reg[10][5]  ( .D(n562), .C(CLK), .Q(\x[10][5] ) );
  DF3 \x_reg[10][4]  ( .D(n561), .C(CLK), .Q(\x[10][4] ) );
  DF3 \x_reg[10][3]  ( .D(n560), .C(CLK), .Q(\x[10][3] ) );
  DF3 \x_reg[10][2]  ( .D(n559), .C(CLK), .Q(\x[10][2] ) );
  DF3 \x_reg[10][1]  ( .D(n558), .C(CLK), .Q(\x[10][1] ) );
  DF3 \x_reg[10][0]  ( .D(n557), .C(CLK), .Q(\x[10][0] ) );
  DF3 \x_reg[11][7]  ( .D(n556), .C(CLK), .Q(\x[11][7] ) );
  DF3 \x_reg[11][6]  ( .D(n555), .C(CLK), .Q(\x[11][6] ) );
  DF3 \x_reg[11][5]  ( .D(n554), .C(CLK), .Q(\x[11][5] ) );
  DF3 \x_reg[11][4]  ( .D(n553), .C(CLK), .Q(\x[11][4] ) );
  DF3 \x_reg[11][3]  ( .D(n552), .C(CLK), .Q(\x[11][3] ) );
  DF3 \x_reg[11][2]  ( .D(n551), .C(CLK), .Q(\x[11][2] ) );
  DF3 \x_reg[11][1]  ( .D(n550), .C(CLK), .Q(\x[11][1] ) );
  DF3 \x_reg[11][0]  ( .D(n549), .C(CLK), .Q(\x[11][0] ) );
  DF3 \x_reg[12][7]  ( .D(n548), .C(CLK), .Q(\x[12][7] ) );
  DF3 \x_reg[12][6]  ( .D(n547), .C(CLK), .Q(\x[12][6] ) );
  DF3 \x_reg[12][5]  ( .D(n546), .C(CLK), .Q(\x[12][5] ) );
  DF3 \x_reg[12][4]  ( .D(n545), .C(CLK), .Q(\x[12][4] ) );
  DF3 \x_reg[12][3]  ( .D(n544), .C(CLK), .Q(\x[12][3] ) );
  DF3 \x_reg[12][2]  ( .D(n543), .C(CLK), .Q(\x[12][2] ) );
  DF3 \x_reg[12][1]  ( .D(n542), .C(CLK), .Q(\x[12][1] ) );
  DF3 \x_reg[12][0]  ( .D(n541), .C(CLK), .Q(\x[12][0] ) );
  DF3 \x_reg[13][7]  ( .D(n540), .C(CLK), .Q(\x[13][7] ) );
  DF3 \x_reg[13][6]  ( .D(n539), .C(CLK), .Q(\x[13][6] ) );
  DF3 \x_reg[13][5]  ( .D(n538), .C(CLK), .Q(\x[13][5] ) );
  DF3 \x_reg[13][4]  ( .D(n537), .C(CLK), .Q(\x[13][4] ) );
  DF3 \x_reg[13][3]  ( .D(n536), .C(CLK), .Q(\x[13][3] ) );
  DF3 \x_reg[13][2]  ( .D(n535), .C(CLK), .Q(\x[13][2] ) );
  DF3 \x_reg[13][1]  ( .D(n534), .C(CLK), .Q(\x[13][1] ) );
  DF3 \x_reg[13][0]  ( .D(n533), .C(CLK), .Q(\x[13][0] ) );
  DF3 \x_reg[14][7]  ( .D(n532), .C(CLK), .Q(\x[14][7] ) );
  DF3 \x_reg[14][6]  ( .D(n531), .C(CLK), .Q(\x[14][6] ) );
  DF3 \x_reg[14][5]  ( .D(n530), .C(CLK), .Q(\x[14][5] ) );
  DF3 \x_reg[14][4]  ( .D(n529), .C(CLK), .Q(\x[14][4] ) );
  DF3 \x_reg[14][3]  ( .D(n528), .C(CLK), .Q(\x[14][3] ) );
  DF3 \x_reg[14][2]  ( .D(n527), .C(CLK), .Q(\x[14][2] ) );
  DF3 \x_reg[14][1]  ( .D(n526), .C(CLK), .Q(\x[14][1] ) );
  DF3 \x_reg[14][0]  ( .D(n525), .C(CLK), .Q(\x[14][0] ) );
  DF3 \x_reg[15][7]  ( .D(n524), .C(CLK), .Q(\x[15][7] ) );
  DF3 \x_reg[15][6]  ( .D(n257), .C(CLK), .Q(\x[15][6] ) );
  DF3 \x_reg[15][5]  ( .D(n248), .C(CLK), .Q(\x[15][5] ) );
  DF3 \x_reg[15][4]  ( .D(n247), .C(CLK), .Q(\x[15][4] ) );
  DF3 \x_reg[15][3]  ( .D(n246), .C(CLK), .Q(\x[15][3] ) );
  DF3 \x_reg[15][2]  ( .D(n245), .C(CLK), .Q(\x[15][2] ) );
  DF3 \x_reg[15][1]  ( .D(n244), .C(CLK), .Q(\x[15][1] ) );
  DF3 \x_reg[15][0]  ( .D(n243), .C(CLK), .Q(\x[15][0] ) );
  DF3 \x_reg[16][7]  ( .D(n242), .C(CLK), .Q(\x[16][7] ) );
  DF3 \x_reg[16][6]  ( .D(n241), .C(CLK), .Q(\x[16][6] ) );
  DF3 \x_reg[16][5]  ( .D(n240), .C(CLK), .Q(\x[16][5] ) );
  DF3 \x_reg[16][4]  ( .D(n239), .C(CLK), .Q(\x[16][4] ) );
  DF3 \x_reg[16][3]  ( .D(n238), .C(CLK), .Q(\x[16][3] ) );
  DF3 \x_reg[16][2]  ( .D(n237), .C(CLK), .Q(\x[16][2] ) );
  DF3 \x_reg[16][1]  ( .D(n236), .C(CLK), .Q(\x[16][1] ) );
  DF3 \x_reg[16][0]  ( .D(n235), .C(CLK), .Q(\x[16][0] ) );
  DF3 \x_reg[17][7]  ( .D(n234), .C(CLK), .Q(\x[17][7] ) );
  DF3 \x_reg[17][6]  ( .D(n233), .C(CLK), .Q(\x[17][6] ) );
  DF3 \x_reg[17][5]  ( .D(n232), .C(CLK), .Q(\x[17][5] ) );
  DF3 \x_reg[17][4]  ( .D(n231), .C(CLK), .Q(\x[17][4] ) );
  DF3 \x_reg[17][3]  ( .D(n230), .C(CLK), .Q(\x[17][3] ) );
  DF3 \x_reg[17][2]  ( .D(n229), .C(CLK), .Q(\x[17][2] ) );
  DF3 \x_reg[17][1]  ( .D(n228), .C(CLK), .Q(\x[17][1] ) );
  DF3 \x_reg[17][0]  ( .D(n227), .C(CLK), .Q(\x[17][0] ) );
  DF3 \x_reg[18][7]  ( .D(n226), .C(CLK), .Q(\x[18][7] ) );
  DF3 \x_reg[18][6]  ( .D(n225), .C(CLK), .Q(\x[18][6] ) );
  DF3 \x_reg[18][5]  ( .D(n224), .C(CLK), .Q(\x[18][5] ) );
  DF3 \x_reg[18][4]  ( .D(n223), .C(CLK), .Q(\x[18][4] ) );
  DF3 \x_reg[18][3]  ( .D(n222), .C(CLK), .Q(\x[18][3] ) );
  DF3 \x_reg[18][2]  ( .D(n221), .C(CLK), .Q(\x[18][2] ) );
  DF3 \x_reg[18][1]  ( .D(n220), .C(CLK), .Q(\x[18][1] ) );
  DF3 \x_reg[18][0]  ( .D(n219), .C(CLK), .Q(\x[18][0] ) );
  DF3 \x_reg[19][7]  ( .D(n218), .C(CLK), .Q(\x[19][7] ) );
  DF3 \x_reg[19][6]  ( .D(n217), .C(CLK), .Q(\x[19][6] ) );
  DF3 \x_reg[19][5]  ( .D(n216), .C(CLK), .Q(\x[19][5] ) );
  DF3 \x_reg[19][4]  ( .D(n215), .C(CLK), .Q(\x[19][4] ) );
  DF3 \x_reg[19][3]  ( .D(n214), .C(CLK), .Q(\x[19][3] ) );
  DF3 \x_reg[19][2]  ( .D(n213), .C(CLK), .Q(\x[19][2] ) );
  DF3 \x_reg[19][1]  ( .D(n212), .C(CLK), .Q(\x[19][1] ) );
  DF3 \x_reg[19][0]  ( .D(n211), .C(CLK), .Q(\x[19][0] ) );
  DF3 \x_reg[20][7]  ( .D(n210), .C(CLK), .Q(\x[20][7] ) );
  DF3 \x_reg[20][6]  ( .D(n209), .C(CLK), .Q(\x[20][6] ) );
  DF3 \x_reg[20][5]  ( .D(n208), .C(CLK), .Q(\x[20][5] ) );
  DF3 \x_reg[20][4]  ( .D(n207), .C(CLK), .Q(\x[20][4] ) );
  DF3 \x_reg[20][3]  ( .D(n206), .C(CLK), .Q(\x[20][3] ) );
  DF3 \x_reg[20][2]  ( .D(n205), .C(CLK), .Q(\x[20][2] ) );
  DF3 \x_reg[20][1]  ( .D(n204), .C(CLK), .Q(\x[20][1] ) );
  DF3 \x_reg[20][0]  ( .D(n203), .C(CLK), .Q(\x[20][0] ) );
  DF3 \x_reg[21][7]  ( .D(n202), .C(CLK), .Q(\x[21][7] ) );
  DF3 \x_reg[21][6]  ( .D(n201), .C(CLK), .Q(\x[21][6] ) );
  DF3 \x_reg[21][5]  ( .D(n200), .C(CLK), .Q(\x[21][5] ) );
  DF3 \x_reg[21][4]  ( .D(n199), .C(CLK), .Q(\x[21][4] ) );
  DF3 \x_reg[21][3]  ( .D(n198), .C(CLK), .Q(\x[21][3] ) );
  DF3 \x_reg[21][2]  ( .D(n197), .C(CLK), .Q(\x[21][2] ) );
  DF3 \x_reg[21][1]  ( .D(n196), .C(CLK), .Q(\x[21][1] ) );
  DF3 \x_reg[21][0]  ( .D(n195), .C(CLK), .Q(\x[21][0] ) );
  DF3 \x_reg[22][7]  ( .D(n194), .C(CLK), .Q(\x[22][7] ) );
  DF3 \x_reg[22][6]  ( .D(n193), .C(CLK), .Q(\x[22][6] ) );
  DF3 \x_reg[22][5]  ( .D(n192), .C(CLK), .Q(\x[22][5] ) );
  DF3 \x_reg[22][4]  ( .D(n191), .C(CLK), .Q(\x[22][4] ) );
  DF3 \x_reg[22][3]  ( .D(n190), .C(CLK), .Q(\x[22][3] ) );
  DF3 \x_reg[22][2]  ( .D(n189), .C(CLK), .Q(\x[22][2] ) );
  DF3 \x_reg[22][1]  ( .D(n188), .C(CLK), .Q(\x[22][1] ) );
  DF3 \x_reg[22][0]  ( .D(n187), .C(CLK), .Q(\x[22][0] ) );
  DF3 \x_reg[23][7]  ( .D(n186), .C(CLK), .Q(\x[23][7] ) );
  DF3 \x_reg[23][6]  ( .D(n185), .C(CLK), .Q(\x[23][6] ) );
  DF3 \x_reg[23][5]  ( .D(n184), .C(CLK), .Q(\x[23][5] ) );
  DF3 \x_reg[23][4]  ( .D(n183), .C(CLK), .Q(\x[23][4] ) );
  DF3 \x_reg[23][3]  ( .D(n182), .C(CLK), .Q(\x[23][3] ) );
  DF3 \x_reg[23][2]  ( .D(n181), .C(CLK), .Q(\x[23][2] ) );
  DF3 \x_reg[23][1]  ( .D(n180), .C(CLK), .Q(\x[23][1] ) );
  DF3 \x_reg[23][0]  ( .D(n179), .C(CLK), .Q(\x[23][0] ) );
  DF3 \x_reg[24][7]  ( .D(n178), .C(CLK), .Q(\x[24][7] ) );
  DF3 \x_reg[24][6]  ( .D(n177), .C(CLK), .Q(\x[24][6] ) );
  DF3 \x_reg[24][5]  ( .D(n176), .C(CLK), .Q(\x[24][5] ) );
  DF3 \x_reg[24][4]  ( .D(n175), .C(CLK), .Q(\x[24][4] ) );
  DF3 \x_reg[24][3]  ( .D(n174), .C(CLK), .Q(\x[24][3] ) );
  DF3 \x_reg[24][2]  ( .D(n173), .C(CLK), .Q(\x[24][2] ) );
  DF3 \x_reg[24][1]  ( .D(n172), .C(CLK), .Q(\x[24][1] ) );
  DF3 \x_reg[24][0]  ( .D(n171), .C(CLK), .Q(\x[24][0] ) );
  DF3 \x_reg[25][7]  ( .D(n170), .C(CLK), .Q(\x[25][7] ) );
  DF3 \x_reg[25][6]  ( .D(n169), .C(CLK), .Q(\x[25][6] ) );
  DF3 \x_reg[25][5]  ( .D(n168), .C(CLK), .Q(\x[25][5] ) );
  DF3 \x_reg[25][4]  ( .D(n167), .C(CLK), .Q(\x[25][4] ) );
  DF3 \x_reg[25][3]  ( .D(n166), .C(CLK), .Q(\x[25][3] ) );
  DF3 \x_reg[25][2]  ( .D(n165), .C(CLK), .Q(\x[25][2] ) );
  DF3 \x_reg[25][1]  ( .D(n164), .C(CLK), .Q(\x[25][1] ) );
  DF3 \x_reg[25][0]  ( .D(n163), .C(CLK), .Q(\x[25][0] ) );
  DF3 \x_reg[26][7]  ( .D(n162), .C(CLK), .Q(\x[26][7] ) );
  DF3 \x_reg[26][6]  ( .D(n161), .C(CLK), .Q(\x[26][6] ) );
  DF3 \x_reg[26][5]  ( .D(n160), .C(CLK), .Q(\x[26][5] ) );
  DF3 \x_reg[26][4]  ( .D(n159), .C(CLK), .Q(\x[26][4] ) );
  DF3 \x_reg[26][3]  ( .D(n158), .C(CLK), .Q(\x[26][3] ) );
  DF3 \x_reg[26][2]  ( .D(n157), .C(CLK), .Q(\x[26][2] ) );
  DF3 \x_reg[26][1]  ( .D(n156), .C(CLK), .Q(\x[26][1] ) );
  DF3 \x_reg[26][0]  ( .D(n155), .C(CLK), .Q(\x[26][0] ) );
  DF3 \x_reg[27][7]  ( .D(n154), .C(CLK), .Q(\x[27][7] ) );
  DF3 \x_reg[27][6]  ( .D(n153), .C(CLK), .Q(\x[27][6] ) );
  DF3 \x_reg[27][5]  ( .D(n152), .C(CLK), .Q(\x[27][5] ) );
  DF3 \x_reg[27][4]  ( .D(n151), .C(CLK), .Q(\x[27][4] ) );
  DF3 \x_reg[27][3]  ( .D(n150), .C(CLK), .Q(\x[27][3] ) );
  DF3 \x_reg[27][2]  ( .D(n149), .C(CLK), .Q(\x[27][2] ) );
  DF3 \x_reg[27][1]  ( .D(n148), .C(CLK), .Q(\x[27][1] ) );
  DF3 \x_reg[27][0]  ( .D(n147), .C(CLK), .Q(\x[27][0] ) );
  DF3 \x_reg[28][7]  ( .D(n146), .C(CLK), .Q(\x[28][7] ) );
  DF3 \x_reg[28][6]  ( .D(n145), .C(CLK), .Q(\x[28][6] ) );
  DF3 \x_reg[28][5]  ( .D(n144), .C(CLK), .Q(\x[28][5] ) );
  DF3 \x_reg[28][4]  ( .D(n143), .C(CLK), .Q(\x[28][4] ) );
  DF3 \x_reg[28][3]  ( .D(n142), .C(CLK), .Q(\x[28][3] ) );
  DF3 \x_reg[28][2]  ( .D(n141), .C(CLK), .Q(\x[28][2] ) );
  DF3 \x_reg[28][1]  ( .D(n140), .C(CLK), .Q(\x[28][1] ) );
  DF3 \x_reg[28][0]  ( .D(n139), .C(CLK), .Q(\x[28][0] ) );
  DF3 \x_reg[29][7]  ( .D(n138), .C(CLK), .Q(\x[29][7] ) );
  DF3 \x_reg[29][6]  ( .D(n137), .C(CLK), .Q(\x[29][6] ) );
  DF3 \x_reg[29][5]  ( .D(n136), .C(CLK), .Q(\x[29][5] ) );
  DF3 \x_reg[29][4]  ( .D(n135), .C(CLK), .Q(\x[29][4] ) );
  DF3 \x_reg[29][3]  ( .D(n134), .C(CLK), .Q(\x[29][3] ) );
  DF3 \x_reg[29][2]  ( .D(n133), .C(CLK), .Q(\x[29][2] ) );
  DF3 \x_reg[29][1]  ( .D(n132), .C(CLK), .Q(\x[29][1] ) );
  DF3 \x_reg[29][0]  ( .D(n131), .C(CLK), .Q(\x[29][0] ) );
  DF3 \x_reg[30][7]  ( .D(n130), .C(CLK), .Q(\x[30][7] ), .QN(n249) );
  DF3 \x_reg[30][6]  ( .D(n129), .C(CLK), .Q(\x[30][6] ), .QN(n250) );
  DF3 \x_reg[30][5]  ( .D(n128), .C(CLK), .Q(\x[30][5] ), .QN(n251) );
  DF3 \x_reg[30][4]  ( .D(n127), .C(CLK), .Q(\x[30][4] ), .QN(n252) );
  DF3 \x_reg[30][3]  ( .D(n126), .C(CLK), .Q(\x[30][3] ), .QN(n253) );
  DF3 \x_reg[30][2]  ( .D(n125), .C(CLK), .Q(\x[30][2] ), .QN(n254) );
  DF3 \x_reg[30][1]  ( .D(n124), .C(CLK), .Q(\x[30][1] ), .QN(n255) );
  DF3 \x_reg[30][0]  ( .D(n123), .C(CLK), .Q(\x[30][0] ), .QN(n256) );
  DF3 \x_reg[31][7]  ( .D(n523), .C(CLK), .Q(\x[31][7] ) );
  DF3 \x_reg[31][6]  ( .D(n522), .C(CLK), .Q(\x[31][6] ) );
  DF3 \x_reg[31][5]  ( .D(n521), .C(CLK), .Q(\x[31][5] ) );
  DF3 \x_reg[31][4]  ( .D(n520), .C(CLK), .Q(\x[31][4] ) );
  DF3 \x_reg[31][3]  ( .D(n519), .C(CLK), .Q(\x[31][3] ) );
  DF3 \x_reg[31][2]  ( .D(n518), .C(CLK), .Q(\x[31][2] ) );
  DF3 \x_reg[31][1]  ( .D(n517), .C(CLK), .Q(\x[31][1] ) );
  DF3 \x_reg[31][0]  ( .D(n516), .C(CLK), .Q(\x[31][0] ) );
  NOR21 U4 ( .A(n114), .B(RESET), .Q(n267) );
  BUF2 U6 ( .A(N2), .Q(n92) );
  BUF2 U8 ( .A(N2), .Q(n91) );
  BUF2 U10 ( .A(N2), .Q(n93) );
  BUF2 U12 ( .A(n95), .Q(n114) );
  INV3 U14 ( .A(n113), .Q(n96) );
  INV3 U16 ( .A(n111), .Q(n110) );
  INV3 U18 ( .A(n111), .Q(n109) );
  INV3 U19 ( .A(n112), .Q(n108) );
  INV3 U20 ( .A(n112), .Q(n107) );
  INV3 U21 ( .A(n112), .Q(n106) );
  INV3 U22 ( .A(n112), .Q(n105) );
  INV3 U23 ( .A(n112), .Q(n104) );
  INV3 U24 ( .A(n111), .Q(n103) );
  INV3 U25 ( .A(n111), .Q(n102) );
  INV3 U26 ( .A(n112), .Q(n101) );
  INV3 U27 ( .A(n113), .Q(n100) );
  INV3 U28 ( .A(n111), .Q(n99) );
  INV3 U29 ( .A(n112), .Q(n98) );
  INV3 U30 ( .A(n112), .Q(n97) );
  BUF2 U31 ( .A(n95), .Q(n118) );
  BUF2 U32 ( .A(n95), .Q(n120) );
  BUF2 U33 ( .A(n95), .Q(n115) );
  BUF2 U34 ( .A(n122), .Q(n117) );
  BUF2 U35 ( .A(n122), .Q(n119) );
  BUF2 U36 ( .A(n122), .Q(n121) );
  BUF2 U37 ( .A(n122), .Q(n116) );
  BUF2 U38 ( .A(n95), .Q(n122) );
  BUF2 U39 ( .A(n89), .Q(n84) );
  BUF2 U40 ( .A(n90), .Q(n86) );
  BUF2 U41 ( .A(n89), .Q(n85) );
  BUF2 U42 ( .A(n90), .Q(n87) );
  BUF2 U43 ( .A(n88), .Q(n83) );
  BUF2 U44 ( .A(n88), .Q(n81) );
  BUF2 U45 ( .A(n88), .Q(n82) );
  INV3 U46 ( .A(n267), .Q(n111) );
  INV3 U47 ( .A(n267), .Q(n112) );
  INV3 U48 ( .A(n267), .Q(n113) );
  INV3 U49 ( .A(n94), .Q(n95) );
  IMUX40 U50 ( .A(\x[16][5] ), .B(\x[17][5] ), .C(\x[18][5] ), .D(\x[19][5] ), 
        .S0(n92), .S1(n85), .Q(n52) );
  IMUX40 U51 ( .A(\x[24][5] ), .B(\x[25][5] ), .C(\x[26][5] ), .D(\x[27][5] ), 
        .S0(n92), .S1(n85), .Q(n53) );
  IMUX40 U52 ( .A(\x[12][5] ), .B(\x[13][5] ), .C(\x[14][5] ), .D(\x[15][5] ), 
        .S0(n92), .S1(n85), .Q(n60) );
  IMUX40 U53 ( .A(\x[0][5] ), .B(\x[1][5] ), .C(\x[2][5] ), .D(\x[3][5] ), 
        .S0(n92), .S1(n86), .Q(n57) );
  IMUX40 U54 ( .A(\x[8][5] ), .B(\x[9][5] ), .C(\x[10][5] ), .D(\x[11][5] ), 
        .S0(n92), .S1(n85), .Q(n58) );
  IMUX40 U55 ( .A(\x[16][3] ), .B(\x[17][3] ), .C(\x[18][3] ), .D(\x[19][3] ), 
        .S0(n93), .S1(n83), .Q(n32) );
  IMUX40 U56 ( .A(\x[24][3] ), .B(\x[25][3] ), .C(\x[26][3] ), .D(\x[27][3] ), 
        .S0(n91), .S1(n83), .Q(n33) );
  IMUX40 U57 ( .A(\x[12][3] ), .B(\x[13][3] ), .C(\x[14][3] ), .D(\x[15][3] ), 
        .S0(n91), .S1(n84), .Q(n40) );
  IMUX40 U58 ( .A(\x[0][3] ), .B(\x[1][3] ), .C(\x[2][3] ), .D(\x[3][3] ), 
        .S0(n91), .S1(n84), .Q(n37) );
  IMUX40 U59 ( .A(\x[8][3] ), .B(\x[9][3] ), .C(\x[10][3] ), .D(\x[11][3] ), 
        .S0(n91), .S1(n84), .Q(n38) );
  IMUX40 U60 ( .A(\x[16][6] ), .B(\x[17][6] ), .C(\x[18][6] ), .D(\x[19][6] ), 
        .S0(n92), .S1(n86), .Q(n62) );
  IMUX40 U61 ( .A(\x[24][6] ), .B(\x[25][6] ), .C(\x[26][6] ), .D(\x[27][6] ), 
        .S0(n92), .S1(n86), .Q(n63) );
  IMUX40 U62 ( .A(\x[12][6] ), .B(\x[13][6] ), .C(\x[14][6] ), .D(\x[15][6] ), 
        .S0(n93), .S1(n86), .Q(n70) );
  IMUX40 U63 ( .A(\x[0][6] ), .B(\x[1][6] ), .C(\x[2][6] ), .D(\x[3][6] ), 
        .S0(n93), .S1(n87), .Q(n67) );
  IMUX40 U64 ( .A(\x[8][6] ), .B(\x[9][6] ), .C(\x[10][6] ), .D(\x[11][6] ), 
        .S0(n93), .S1(n86), .Q(n68) );
  IMUX40 U65 ( .A(\x[16][4] ), .B(\x[17][4] ), .C(\x[18][4] ), .D(\x[19][4] ), 
        .S0(n91), .S1(n84), .Q(n42) );
  IMUX40 U66 ( .A(\x[24][4] ), .B(\x[25][4] ), .C(\x[26][4] ), .D(\x[27][4] ), 
        .S0(n91), .S1(n84), .Q(n43) );
  IMUX40 U67 ( .A(\x[12][4] ), .B(\x[13][4] ), .C(\x[14][4] ), .D(\x[15][4] ), 
        .S0(n91), .S1(n84), .Q(n50) );
  IMUX40 U68 ( .A(\x[0][4] ), .B(\x[1][4] ), .C(\x[2][4] ), .D(\x[3][4] ), 
        .S0(n91), .S1(n85), .Q(n47) );
  IMUX40 U69 ( .A(\x[8][4] ), .B(\x[9][4] ), .C(\x[10][4] ), .D(\x[11][4] ), 
        .S0(n91), .S1(n85), .Q(n48) );
  IMUX40 U70 ( .A(\x[16][7] ), .B(\x[17][7] ), .C(\x[18][7] ), .D(\x[19][7] ), 
        .S0(n93), .S1(n87), .Q(n72) );
  IMUX40 U71 ( .A(\x[24][7] ), .B(\x[25][7] ), .C(\x[26][7] ), .D(\x[27][7] ), 
        .S0(n93), .S1(n87), .Q(n73) );
  IMUX40 U72 ( .A(\x[12][7] ), .B(\x[13][7] ), .C(\x[14][7] ), .D(\x[15][7] ), 
        .S0(n93), .S1(n87), .Q(n80) );
  IMUX40 U73 ( .A(\x[0][7] ), .B(\x[1][7] ), .C(\x[2][7] ), .D(\x[3][7] ), 
        .S0(n93), .S1(n87), .Q(n77) );
  IMUX40 U74 ( .A(\x[8][7] ), .B(\x[9][7] ), .C(\x[10][7] ), .D(\x[11][7] ), 
        .S0(n93), .S1(n87), .Q(n78) );
  IMUX40 U75 ( .A(\x[28][5] ), .B(\x[29][5] ), .C(\x[30][5] ), .D(\x[31][5] ), 
        .S0(n92), .S1(n85), .Q(n55) );
  IMUX40 U76 ( .A(\x[28][3] ), .B(\x[29][3] ), .C(\x[30][3] ), .D(\x[31][3] ), 
        .S0(n91), .S1(n83), .Q(n35) );
  IMUX40 U77 ( .A(\x[28][6] ), .B(\x[29][6] ), .C(\x[30][6] ), .D(\x[31][6] ), 
        .S0(n92), .S1(n86), .Q(n65) );
  IMUX40 U78 ( .A(\x[28][4] ), .B(\x[29][4] ), .C(\x[30][4] ), .D(\x[31][4] ), 
        .S0(n91), .S1(n84), .Q(n45) );
  IMUX40 U79 ( .A(\x[28][7] ), .B(\x[29][7] ), .C(\x[30][7] ), .D(\x[31][7] ), 
        .S0(n93), .S1(n87), .Q(n75) );
  IMUX40 U80 ( .A(\x[20][5] ), .B(\x[21][5] ), .C(\x[22][5] ), .D(\x[23][5] ), 
        .S0(n92), .S1(n85), .Q(n54) );
  IMUX40 U81 ( .A(\x[20][3] ), .B(\x[21][3] ), .C(\x[22][3] ), .D(\x[23][3] ), 
        .S0(n91), .S1(n83), .Q(n34) );
  IMUX40 U82 ( .A(\x[20][6] ), .B(\x[21][6] ), .C(\x[22][6] ), .D(\x[23][6] ), 
        .S0(n92), .S1(n86), .Q(n64) );
  IMUX40 U83 ( .A(\x[20][4] ), .B(\x[21][4] ), .C(\x[22][4] ), .D(\x[23][4] ), 
        .S0(n91), .S1(n84), .Q(n44) );
  IMUX40 U84 ( .A(\x[20][7] ), .B(\x[21][7] ), .C(\x[22][7] ), .D(\x[23][7] ), 
        .S0(n93), .S1(n87), .Q(n74) );
  MUX22 U85 ( .A(n76), .B(n71), .S(N6), .Q(Delay_Line_out[7]) );
  IMUX40 U86 ( .A(n77), .B(n78), .C(n79), .D(n80), .S0(N5), .S1(N4), .Q(n76)
         );
  IMUX40 U87 ( .A(n72), .B(n73), .C(n74), .D(n75), .S0(N5), .S1(N4), .Q(n71)
         );
  IMUX40 U88 ( .A(\x[4][7] ), .B(\x[5][7] ), .C(\x[6][7] ), .D(\x[7][7] ), 
        .S0(n93), .S1(n87), .Q(n79) );
  MUX22 U89 ( .A(n56), .B(n51), .S(N6), .Q(Delay_Line_out[5]) );
  IMUX40 U90 ( .A(n57), .B(n58), .C(n59), .D(n60), .S0(N5), .S1(N4), .Q(n56)
         );
  IMUX40 U91 ( .A(n52), .B(n53), .C(n54), .D(n55), .S0(N5), .S1(N4), .Q(n51)
         );
  IMUX40 U92 ( .A(\x[4][5] ), .B(\x[5][5] ), .C(\x[6][5] ), .D(\x[7][5] ), 
        .S0(n92), .S1(n86), .Q(n59) );
  MUX22 U93 ( .A(n36), .B(n31), .S(N6), .Q(Delay_Line_out[3]) );
  IMUX40 U94 ( .A(n37), .B(n38), .C(n39), .D(n40), .S0(N5), .S1(N4), .Q(n36)
         );
  IMUX40 U95 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(N5), .S1(N4), .Q(n31)
         );
  IMUX40 U96 ( .A(\x[4][3] ), .B(\x[5][3] ), .C(\x[6][3] ), .D(\x[7][3] ), 
        .S0(n91), .S1(n84), .Q(n39) );
  MUX22 U97 ( .A(n66), .B(n61), .S(N6), .Q(Delay_Line_out[6]) );
  IMUX40 U98 ( .A(n67), .B(n68), .C(n69), .D(n70), .S0(N5), .S1(N4), .Q(n66)
         );
  IMUX40 U99 ( .A(n62), .B(n63), .C(n64), .D(n65), .S0(N5), .S1(N4), .Q(n61)
         );
  IMUX40 U100 ( .A(\x[4][6] ), .B(\x[5][6] ), .C(\x[6][6] ), .D(\x[7][6] ), 
        .S0(n93), .S1(n86), .Q(n69) );
  MUX22 U101 ( .A(n46), .B(n41), .S(N6), .Q(Delay_Line_out[4]) );
  IMUX40 U102 ( .A(n47), .B(n48), .C(n49), .D(n50), .S0(N5), .S1(N4), .Q(n46)
         );
  IMUX40 U103 ( .A(n42), .B(n43), .C(n44), .D(n45), .S0(N5), .S1(N4), .Q(n41)
         );
  IMUX40 U104 ( .A(\x[4][4] ), .B(\x[5][4] ), .C(\x[6][4] ), .D(\x[7][4] ), 
        .S0(n91), .S1(n85), .Q(n49) );
  BUF2 U105 ( .A(N3), .Q(n89) );
  BUF2 U106 ( .A(N3), .Q(n90) );
  IMUX40 U107 ( .A(\x[16][2] ), .B(\x[17][2] ), .C(\x[18][2] ), .D(\x[19][2] ), 
        .S0(n92), .S1(n83), .Q(n22) );
  IMUX40 U108 ( .A(\x[24][2] ), .B(\x[25][2] ), .C(\x[26][2] ), .D(\x[27][2] ), 
        .S0(n92), .S1(n82), .Q(n23) );
  IMUX40 U109 ( .A(\x[12][2] ), .B(\x[13][2] ), .C(\x[14][2] ), .D(\x[15][2] ), 
        .S0(n91), .S1(n83), .Q(n30) );
  IMUX40 U110 ( .A(\x[8][2] ), .B(\x[9][2] ), .C(\x[10][2] ), .D(\x[11][2] ), 
        .S0(n91), .S1(n83), .Q(n28) );
  IMUX40 U111 ( .A(\x[0][2] ), .B(\x[1][2] ), .C(\x[2][2] ), .D(\x[3][2] ), 
        .S0(n91), .S1(n83), .Q(n27) );
  IMUX40 U112 ( .A(\x[12][0] ), .B(\x[13][0] ), .C(\x[14][0] ), .D(\x[15][0] ), 
        .S0(N2), .S1(n81), .Q(n10) );
  IMUX40 U113 ( .A(\x[0][0] ), .B(\x[1][0] ), .C(\x[2][0] ), .D(\x[3][0] ), 
        .S0(N2), .S1(n81), .Q(n7) );
  IMUX40 U114 ( .A(\x[8][0] ), .B(\x[9][0] ), .C(\x[10][0] ), .D(\x[11][0] ), 
        .S0(N2), .S1(n81), .Q(n8) );
  IMUX40 U115 ( .A(\x[16][0] ), .B(\x[17][0] ), .C(\x[18][0] ), .D(\x[19][0] ), 
        .S0(N2), .S1(n81), .Q(n2) );
  IMUX40 U116 ( .A(\x[24][0] ), .B(\x[25][0] ), .C(\x[26][0] ), .D(\x[27][0] ), 
        .S0(N2), .S1(n81), .Q(n3) );
  IMUX40 U117 ( .A(\x[16][1] ), .B(\x[17][1] ), .C(\x[18][1] ), .D(\x[19][1] ), 
        .S0(N2), .S1(n82), .Q(n12) );
  IMUX40 U118 ( .A(\x[24][1] ), .B(\x[25][1] ), .C(\x[26][1] ), .D(\x[27][1] ), 
        .S0(N2), .S1(n81), .Q(n13) );
  IMUX40 U119 ( .A(\x[12][1] ), .B(\x[13][1] ), .C(\x[14][1] ), .D(\x[15][1] ), 
        .S0(n93), .S1(n82), .Q(n20) );
  IMUX40 U120 ( .A(\x[8][1] ), .B(\x[9][1] ), .C(\x[10][1] ), .D(\x[11][1] ), 
        .S0(N2), .S1(n82), .Q(n18) );
  IMUX40 U121 ( .A(\x[0][1] ), .B(\x[1][1] ), .C(\x[2][1] ), .D(\x[3][1] ), 
        .S0(N2), .S1(n82), .Q(n17) );
  IMUX40 U122 ( .A(\x[28][2] ), .B(\x[29][2] ), .C(\x[30][2] ), .D(\x[31][2] ), 
        .S0(n92), .S1(n82), .Q(n25) );
  IMUX40 U123 ( .A(\x[28][1] ), .B(\x[29][1] ), .C(\x[30][1] ), .D(\x[31][1] ), 
        .S0(N2), .S1(n81), .Q(n15) );
  IMUX40 U124 ( .A(\x[20][2] ), .B(\x[21][2] ), .C(\x[22][2] ), .D(\x[23][2] ), 
        .S0(n93), .S1(n82), .Q(n24) );
  IMUX40 U125 ( .A(\x[4][0] ), .B(\x[5][0] ), .C(\x[6][0] ), .D(\x[7][0] ), 
        .S0(N2), .S1(n81), .Q(n9) );
  IMUX40 U126 ( .A(\x[20][0] ), .B(\x[21][0] ), .C(\x[22][0] ), .D(\x[23][0] ), 
        .S0(N2), .S1(n81), .Q(n4) );
  IMUX40 U127 ( .A(\x[20][1] ), .B(\x[21][1] ), .C(\x[22][1] ), .D(\x[23][1] ), 
        .S0(N2), .S1(n82), .Q(n14) );
  MUX22 U128 ( .A(n26), .B(n21), .S(N6), .Q(Delay_Line_out[2]) );
  IMUX40 U129 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(N5), .S1(N4), .Q(n26)
         );
  IMUX40 U130 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(N5), .S1(N4), .Q(n21)
         );
  IMUX40 U131 ( .A(\x[4][2] ), .B(\x[5][2] ), .C(\x[6][2] ), .D(\x[7][2] ), 
        .S0(n92), .S1(n83), .Q(n29) );
  MUX22 U132 ( .A(n6), .B(n1), .S(N6), .Q(Delay_Line_out[0]) );
  IMUX40 U133 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(N5), .S1(N4), .Q(n1) );
  IMUX40 U134 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(N5), .S1(N4), .Q(n6) );
  IMUX40 U135 ( .A(\x[28][0] ), .B(\x[29][0] ), .C(\x[30][0] ), .D(\x[31][0] ), 
        .S0(N2), .S1(n81), .Q(n5) );
  MUX22 U136 ( .A(n16), .B(n11), .S(N6), .Q(Delay_Line_out[1]) );
  IMUX40 U137 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(N5), .S1(N4), .Q(n16)
         );
  IMUX40 U138 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(N5), .S1(N4), .Q(n11)
         );
  IMUX40 U139 ( .A(\x[4][1] ), .B(\x[5][1] ), .C(\x[6][1] ), .D(\x[7][1] ), 
        .S0(N2), .S1(n82), .Q(n19) );
  BUF2 U140 ( .A(N3), .Q(n88) );
  INV3 U141 ( .A(n387), .Q(n525) );
  AOI221 U142 ( .A(n122), .B(\x[14][0] ), .C(n103), .D(\x[13][0] ), .Q(n387)
         );
  INV3 U143 ( .A(n388), .Q(n524) );
  AOI221 U144 ( .A(n122), .B(\x[15][7] ), .C(n103), .D(\x[14][7] ), .Q(n388)
         );
  NAND22 U145 ( .A(\x[31][3] ), .B(n114), .Q(n262) );
  NAND22 U146 ( .A(\x[31][4] ), .B(n114), .Q(n263) );
  NAND22 U147 ( .A(\x[31][5] ), .B(n114), .Q(n264) );
  NAND22 U148 ( .A(\x[31][6] ), .B(n114), .Q(n265) );
  NAND22 U149 ( .A(\x[31][7] ), .B(n114), .Q(n266) );
  INV3 U150 ( .A(n259), .Q(n94) );
  NOR21 U151 ( .A(RESET), .B(Delay_Line_sample_shift), .Q(n259) );
  INV3 U152 ( .A(n512), .Q(n126) );
  AOI221 U153 ( .A(n118), .B(\x[30][3] ), .C(n103), .D(\x[29][3] ), .Q(n512)
         );
  INV3 U154 ( .A(n511), .Q(n127) );
  AOI221 U155 ( .A(n120), .B(\x[30][4] ), .C(n99), .D(\x[29][4] ), .Q(n511) );
  INV3 U156 ( .A(n510), .Q(n128) );
  AOI221 U157 ( .A(n115), .B(\x[30][5] ), .C(n102), .D(\x[29][5] ), .Q(n510)
         );
  INV3 U158 ( .A(n509), .Q(n129) );
  AOI221 U159 ( .A(n115), .B(\x[30][6] ), .C(n110), .D(\x[29][6] ), .Q(n509)
         );
  INV3 U160 ( .A(n508), .Q(n130) );
  AOI221 U161 ( .A(n118), .B(\x[30][7] ), .C(n109), .D(\x[29][7] ), .Q(n508)
         );
  INV3 U162 ( .A(n507), .Q(n131) );
  AOI221 U163 ( .A(n120), .B(\x[29][0] ), .C(n103), .D(\x[28][0] ), .Q(n507)
         );
  INV3 U164 ( .A(n506), .Q(n132) );
  AOI221 U165 ( .A(n115), .B(\x[29][1] ), .C(n99), .D(\x[28][1] ), .Q(n506) );
  INV3 U166 ( .A(n505), .Q(n133) );
  AOI221 U167 ( .A(n115), .B(\x[29][2] ), .C(n110), .D(\x[28][2] ), .Q(n505)
         );
  INV3 U168 ( .A(n504), .Q(n134) );
  AOI221 U169 ( .A(n118), .B(\x[29][3] ), .C(n110), .D(\x[28][3] ), .Q(n504)
         );
  INV3 U170 ( .A(n503), .Q(n135) );
  AOI221 U171 ( .A(n120), .B(\x[29][4] ), .C(n110), .D(\x[28][4] ), .Q(n503)
         );
  INV3 U172 ( .A(n502), .Q(n136) );
  AOI221 U173 ( .A(n115), .B(\x[29][5] ), .C(n110), .D(\x[28][5] ), .Q(n502)
         );
  INV3 U174 ( .A(n501), .Q(n137) );
  AOI221 U175 ( .A(n118), .B(\x[29][6] ), .C(n110), .D(\x[28][6] ), .Q(n501)
         );
  INV3 U176 ( .A(n500), .Q(n138) );
  AOI221 U177 ( .A(n118), .B(\x[29][7] ), .C(n110), .D(\x[28][7] ), .Q(n500)
         );
  INV3 U178 ( .A(n499), .Q(n139) );
  AOI221 U179 ( .A(n120), .B(\x[28][0] ), .C(n110), .D(\x[27][0] ), .Q(n499)
         );
  INV3 U180 ( .A(n498), .Q(n140) );
  AOI221 U181 ( .A(n115), .B(\x[28][1] ), .C(n110), .D(\x[27][1] ), .Q(n498)
         );
  INV3 U182 ( .A(n475), .Q(n163) );
  AOI221 U183 ( .A(n118), .B(\x[25][0] ), .C(n109), .D(\x[24][0] ), .Q(n475)
         );
  INV3 U184 ( .A(n474), .Q(n164) );
  AOI221 U185 ( .A(n118), .B(\x[25][1] ), .C(n109), .D(\x[24][1] ), .Q(n474)
         );
  INV3 U186 ( .A(n473), .Q(n165) );
  AOI221 U187 ( .A(n118), .B(\x[25][2] ), .C(n108), .D(\x[24][2] ), .Q(n473)
         );
  INV3 U188 ( .A(n472), .Q(n166) );
  AOI221 U189 ( .A(n118), .B(\x[25][3] ), .C(n108), .D(\x[24][3] ), .Q(n472)
         );
  INV3 U190 ( .A(n471), .Q(n167) );
  AOI221 U191 ( .A(n118), .B(\x[25][4] ), .C(n108), .D(\x[24][4] ), .Q(n471)
         );
  INV3 U192 ( .A(n470), .Q(n168) );
  AOI221 U193 ( .A(n118), .B(\x[25][5] ), .C(n108), .D(\x[24][5] ), .Q(n470)
         );
  INV3 U194 ( .A(n469), .Q(n169) );
  AOI221 U195 ( .A(n118), .B(\x[25][6] ), .C(n108), .D(\x[24][6] ), .Q(n469)
         );
  INV3 U196 ( .A(n468), .Q(n170) );
  AOI221 U197 ( .A(n118), .B(\x[25][7] ), .C(n108), .D(\x[24][7] ), .Q(n468)
         );
  INV3 U198 ( .A(n467), .Q(n171) );
  AOI221 U199 ( .A(n118), .B(\x[24][0] ), .C(n108), .D(\x[23][0] ), .Q(n467)
         );
  INV3 U200 ( .A(n466), .Q(n172) );
  AOI221 U201 ( .A(n118), .B(\x[24][1] ), .C(n108), .D(\x[23][1] ), .Q(n466)
         );
  INV3 U202 ( .A(n465), .Q(n173) );
  AOI221 U203 ( .A(n118), .B(\x[24][2] ), .C(n108), .D(\x[23][2] ), .Q(n465)
         );
  INV3 U204 ( .A(n464), .Q(n174) );
  AOI221 U205 ( .A(n118), .B(\x[24][3] ), .C(n108), .D(\x[23][3] ), .Q(n464)
         );
  INV3 U206 ( .A(n463), .Q(n175) );
  AOI221 U207 ( .A(n118), .B(\x[24][4] ), .C(n108), .D(\x[23][4] ), .Q(n463)
         );
  INV3 U208 ( .A(n462), .Q(n176) );
  AOI221 U209 ( .A(n118), .B(\x[24][5] ), .C(n108), .D(\x[23][5] ), .Q(n462)
         );
  INV3 U210 ( .A(n461), .Q(n177) );
  AOI221 U211 ( .A(n118), .B(\x[24][6] ), .C(n108), .D(\x[23][6] ), .Q(n461)
         );
  INV3 U212 ( .A(n460), .Q(n178) );
  AOI221 U213 ( .A(n118), .B(\x[24][7] ), .C(n108), .D(\x[23][7] ), .Q(n460)
         );
  INV3 U214 ( .A(n459), .Q(n179) );
  AOI221 U215 ( .A(n118), .B(\x[23][0] ), .C(n108), .D(\x[22][0] ), .Q(n459)
         );
  INV3 U216 ( .A(n458), .Q(n180) );
  AOI221 U217 ( .A(n118), .B(\x[23][1] ), .C(n108), .D(\x[22][1] ), .Q(n458)
         );
  INV3 U218 ( .A(n457), .Q(n181) );
  AOI221 U219 ( .A(n118), .B(\x[23][2] ), .C(n107), .D(\x[22][2] ), .Q(n457)
         );
  INV3 U220 ( .A(n456), .Q(n182) );
  AOI221 U221 ( .A(n118), .B(\x[23][3] ), .C(n107), .D(\x[22][3] ), .Q(n456)
         );
  INV3 U222 ( .A(n455), .Q(n183) );
  AOI221 U223 ( .A(n118), .B(\x[23][4] ), .C(n107), .D(\x[22][4] ), .Q(n455)
         );
  INV3 U224 ( .A(n454), .Q(n184) );
  AOI221 U225 ( .A(n118), .B(\x[23][5] ), .C(n107), .D(\x[22][5] ), .Q(n454)
         );
  INV3 U226 ( .A(n432), .Q(n206) );
  AOI221 U227 ( .A(n120), .B(\x[20][3] ), .C(n106), .D(\x[19][3] ), .Q(n432)
         );
  INV3 U228 ( .A(n431), .Q(n207) );
  AOI221 U229 ( .A(n120), .B(\x[20][4] ), .C(n106), .D(\x[19][4] ), .Q(n431)
         );
  INV3 U230 ( .A(n430), .Q(n208) );
  AOI221 U231 ( .A(n120), .B(\x[20][5] ), .C(n106), .D(\x[19][5] ), .Q(n430)
         );
  INV3 U232 ( .A(n429), .Q(n209) );
  AOI221 U233 ( .A(n120), .B(\x[20][6] ), .C(n106), .D(\x[19][6] ), .Q(n429)
         );
  INV3 U234 ( .A(n428), .Q(n210) );
  AOI221 U235 ( .A(n120), .B(\x[20][7] ), .C(n106), .D(\x[19][7] ), .Q(n428)
         );
  INV3 U236 ( .A(n427), .Q(n211) );
  AOI221 U237 ( .A(n120), .B(\x[19][0] ), .C(n106), .D(\x[18][0] ), .Q(n427)
         );
  INV3 U238 ( .A(n426), .Q(n212) );
  AOI221 U239 ( .A(n120), .B(\x[19][1] ), .C(n106), .D(\x[18][1] ), .Q(n426)
         );
  INV3 U240 ( .A(n425), .Q(n213) );
  AOI221 U241 ( .A(n120), .B(\x[19][2] ), .C(n105), .D(\x[18][2] ), .Q(n425)
         );
  INV3 U242 ( .A(n424), .Q(n214) );
  AOI221 U243 ( .A(n120), .B(\x[19][3] ), .C(n105), .D(\x[18][3] ), .Q(n424)
         );
  INV3 U244 ( .A(n423), .Q(n215) );
  AOI221 U245 ( .A(n120), .B(\x[19][4] ), .C(n105), .D(\x[18][4] ), .Q(n423)
         );
  INV3 U246 ( .A(n422), .Q(n216) );
  AOI221 U247 ( .A(n120), .B(\x[19][5] ), .C(n105), .D(\x[18][5] ), .Q(n422)
         );
  INV3 U248 ( .A(n421), .Q(n217) );
  AOI221 U249 ( .A(n120), .B(\x[19][6] ), .C(n105), .D(\x[18][6] ), .Q(n421)
         );
  INV3 U250 ( .A(n420), .Q(n218) );
  AOI221 U251 ( .A(n120), .B(\x[19][7] ), .C(n105), .D(\x[18][7] ), .Q(n420)
         );
  INV3 U252 ( .A(n419), .Q(n219) );
  AOI221 U253 ( .A(n120), .B(\x[18][0] ), .C(n105), .D(\x[17][0] ), .Q(n419)
         );
  INV3 U254 ( .A(n418), .Q(n220) );
  AOI221 U255 ( .A(n120), .B(\x[18][1] ), .C(n105), .D(\x[17][1] ), .Q(n418)
         );
  INV3 U256 ( .A(n417), .Q(n221) );
  AOI221 U257 ( .A(n120), .B(\x[18][2] ), .C(n105), .D(\x[17][2] ), .Q(n417)
         );
  INV3 U258 ( .A(n416), .Q(n222) );
  AOI221 U259 ( .A(n120), .B(\x[18][3] ), .C(n105), .D(\x[17][3] ), .Q(n416)
         );
  INV3 U260 ( .A(n415), .Q(n223) );
  AOI221 U261 ( .A(n120), .B(\x[18][4] ), .C(n105), .D(\x[17][4] ), .Q(n415)
         );
  INV3 U262 ( .A(n414), .Q(n224) );
  AOI221 U263 ( .A(n120), .B(\x[18][5] ), .C(n105), .D(\x[17][5] ), .Q(n414)
         );
  INV3 U264 ( .A(n413), .Q(n225) );
  AOI221 U265 ( .A(n120), .B(\x[18][6] ), .C(n105), .D(\x[17][6] ), .Q(n413)
         );
  INV3 U266 ( .A(n412), .Q(n226) );
  AOI221 U267 ( .A(n120), .B(\x[18][7] ), .C(n105), .D(\x[17][7] ), .Q(n412)
         );
  INV3 U268 ( .A(n411), .Q(n227) );
  AOI221 U269 ( .A(n120), .B(\x[17][0] ), .C(n105), .D(\x[16][0] ), .Q(n411)
         );
  INV3 U270 ( .A(n373), .Q(n539) );
  AOI221 U271 ( .A(n115), .B(\x[13][6] ), .C(n102), .D(\x[12][6] ), .Q(n373)
         );
  INV3 U272 ( .A(n368), .Q(n544) );
  AOI221 U273 ( .A(n115), .B(\x[12][3] ), .C(n102), .D(\x[11][3] ), .Q(n368)
         );
  INV3 U274 ( .A(n367), .Q(n545) );
  AOI221 U275 ( .A(n115), .B(\x[12][4] ), .C(n102), .D(\x[11][4] ), .Q(n367)
         );
  INV3 U276 ( .A(n366), .Q(n546) );
  AOI221 U277 ( .A(n115), .B(\x[12][5] ), .C(n102), .D(\x[11][5] ), .Q(n366)
         );
  INV3 U278 ( .A(n365), .Q(n547) );
  AOI221 U279 ( .A(n115), .B(\x[12][6] ), .C(n102), .D(\x[11][6] ), .Q(n365)
         );
  INV3 U280 ( .A(n364), .Q(n548) );
  AOI221 U281 ( .A(n115), .B(\x[12][7] ), .C(n102), .D(\x[11][7] ), .Q(n364)
         );
  INV3 U282 ( .A(n363), .Q(n549) );
  AOI221 U283 ( .A(n115), .B(\x[11][0] ), .C(n102), .D(\x[10][0] ), .Q(n363)
         );
  INV3 U284 ( .A(n362), .Q(n550) );
  AOI221 U285 ( .A(n115), .B(\x[11][1] ), .C(n102), .D(\x[10][1] ), .Q(n362)
         );
  INV3 U286 ( .A(n361), .Q(n551) );
  AOI221 U287 ( .A(n115), .B(\x[11][2] ), .C(n101), .D(\x[10][2] ), .Q(n361)
         );
  INV3 U288 ( .A(n360), .Q(n552) );
  AOI221 U289 ( .A(n115), .B(\x[11][3] ), .C(n101), .D(\x[10][3] ), .Q(n360)
         );
  INV3 U290 ( .A(n359), .Q(n553) );
  AOI221 U291 ( .A(n115), .B(\x[11][4] ), .C(n101), .D(\x[10][4] ), .Q(n359)
         );
  INV3 U292 ( .A(n358), .Q(n554) );
  AOI221 U293 ( .A(n115), .B(\x[11][5] ), .C(n101), .D(\x[10][5] ), .Q(n358)
         );
  INV3 U294 ( .A(n357), .Q(n555) );
  AOI221 U295 ( .A(n115), .B(\x[11][6] ), .C(n101), .D(\x[10][6] ), .Q(n357)
         );
  INV3 U296 ( .A(n356), .Q(n556) );
  AOI221 U297 ( .A(n115), .B(\x[11][7] ), .C(n101), .D(\x[10][7] ), .Q(n356)
         );
  INV3 U298 ( .A(n355), .Q(n557) );
  AOI221 U299 ( .A(n115), .B(\x[10][0] ), .C(n101), .D(\x[9][0] ), .Q(n355) );
  INV3 U300 ( .A(n354), .Q(n558) );
  AOI221 U301 ( .A(n115), .B(\x[10][1] ), .C(n101), .D(\x[9][1] ), .Q(n354) );
  INV3 U302 ( .A(n353), .Q(n559) );
  AOI221 U303 ( .A(n115), .B(\x[10][2] ), .C(n101), .D(\x[9][2] ), .Q(n353) );
  INV3 U304 ( .A(n352), .Q(n560) );
  AOI221 U305 ( .A(n115), .B(\x[10][3] ), .C(n101), .D(\x[9][3] ), .Q(n352) );
  INV3 U306 ( .A(n351), .Q(n561) );
  AOI221 U307 ( .A(n115), .B(\x[10][4] ), .C(n101), .D(\x[9][4] ), .Q(n351) );
  INV3 U308 ( .A(n350), .Q(n562) );
  AOI221 U309 ( .A(n115), .B(\x[10][5] ), .C(n101), .D(\x[9][5] ), .Q(n350) );
  INV3 U310 ( .A(n348), .Q(n564) );
  AOI221 U311 ( .A(n115), .B(\x[10][7] ), .C(n101), .D(\x[9][7] ), .Q(n348) );
  INV3 U312 ( .A(n347), .Q(n565) );
  AOI221 U313 ( .A(n115), .B(\x[9][0] ), .C(n101), .D(\x[8][0] ), .Q(n347) );
  INV3 U314 ( .A(n326), .Q(n586) );
  AOI221 U315 ( .A(n118), .B(\x[7][5] ), .C(n99), .D(\x[6][5] ), .Q(n326) );
  INV3 U316 ( .A(n325), .Q(n587) );
  AOI221 U317 ( .A(n120), .B(\x[7][6] ), .C(n99), .D(\x[6][6] ), .Q(n325) );
  INV3 U318 ( .A(n324), .Q(n588) );
  AOI221 U319 ( .A(n120), .B(\x[7][7] ), .C(n99), .D(\x[6][7] ), .Q(n324) );
  INV3 U320 ( .A(n323), .Q(n589) );
  AOI221 U321 ( .A(n115), .B(\x[6][0] ), .C(n99), .D(\x[5][0] ), .Q(n323) );
  INV3 U322 ( .A(n322), .Q(n590) );
  AOI221 U323 ( .A(n118), .B(\x[6][1] ), .C(n99), .D(\x[5][1] ), .Q(n322) );
  INV3 U324 ( .A(n321), .Q(n591) );
  AOI221 U325 ( .A(n120), .B(\x[6][2] ), .C(n99), .D(\x[5][2] ), .Q(n321) );
  INV3 U326 ( .A(n320), .Q(n592) );
  AOI221 U327 ( .A(n115), .B(\x[6][3] ), .C(n99), .D(\x[5][3] ), .Q(n320) );
  INV3 U328 ( .A(n319), .Q(n593) );
  AOI221 U329 ( .A(n118), .B(\x[6][4] ), .C(n99), .D(\x[5][4] ), .Q(n319) );
  INV3 U330 ( .A(n318), .Q(n594) );
  AOI221 U331 ( .A(n120), .B(\x[6][5] ), .C(n99), .D(\x[5][5] ), .Q(n318) );
  INV3 U332 ( .A(n317), .Q(n595) );
  AOI221 U333 ( .A(n115), .B(\x[6][6] ), .C(n99), .D(\x[5][6] ), .Q(n317) );
  INV3 U334 ( .A(n316), .Q(n596) );
  AOI221 U335 ( .A(n118), .B(\x[6][7] ), .C(n99), .D(\x[5][7] ), .Q(n316) );
  INV3 U336 ( .A(n315), .Q(n597) );
  AOI221 U337 ( .A(n120), .B(\x[5][0] ), .C(n99), .D(\x[4][0] ), .Q(n315) );
  INV3 U338 ( .A(n314), .Q(n598) );
  AOI221 U339 ( .A(n122), .B(\x[5][1] ), .C(n99), .D(\x[4][1] ), .Q(n314) );
  INV3 U340 ( .A(n313), .Q(n599) );
  AOI221 U341 ( .A(n115), .B(\x[5][2] ), .C(n98), .D(\x[4][2] ), .Q(n313) );
  INV3 U342 ( .A(n312), .Q(n600) );
  AOI221 U343 ( .A(n118), .B(\x[5][3] ), .C(n98), .D(\x[4][3] ), .Q(n312) );
  INV3 U344 ( .A(n311), .Q(n601) );
  AOI221 U345 ( .A(n120), .B(\x[5][4] ), .C(n98), .D(\x[4][4] ), .Q(n311) );
  INV3 U346 ( .A(n310), .Q(n602) );
  AOI221 U347 ( .A(n115), .B(\x[5][5] ), .C(n98), .D(\x[4][5] ), .Q(n310) );
  INV3 U348 ( .A(n309), .Q(n603) );
  AOI221 U349 ( .A(n122), .B(\x[5][6] ), .C(n98), .D(\x[4][6] ), .Q(n309) );
  INV3 U350 ( .A(n308), .Q(n604) );
  AOI221 U351 ( .A(n118), .B(\x[5][7] ), .C(n98), .D(\x[4][7] ), .Q(n308) );
  INV3 U352 ( .A(n307), .Q(n605) );
  AOI221 U353 ( .A(n120), .B(\x[4][0] ), .C(n98), .D(\x[3][0] ), .Q(n307) );
  INV3 U354 ( .A(n306), .Q(n606) );
  AOI221 U355 ( .A(n115), .B(\x[4][1] ), .C(n98), .D(\x[3][1] ), .Q(n306) );
  INV3 U356 ( .A(n305), .Q(n607) );
  AOI221 U357 ( .A(n122), .B(\x[4][2] ), .C(n98), .D(\x[3][2] ), .Q(n305) );
  INV3 U358 ( .A(n304), .Q(n608) );
  AOI221 U359 ( .A(n118), .B(\x[4][3] ), .C(n98), .D(\x[3][3] ), .Q(n304) );
  INV3 U360 ( .A(n281), .Q(n631) );
  AOI221 U361 ( .A(n118), .B(\x[1][2] ), .C(n96), .D(\x[0][2] ), .Q(n281) );
  INV3 U362 ( .A(n280), .Q(n632) );
  AOI221 U363 ( .A(n120), .B(\x[1][3] ), .C(n96), .D(\x[0][3] ), .Q(n280) );
  INV3 U364 ( .A(n279), .Q(n633) );
  AOI221 U365 ( .A(n115), .B(\x[1][4] ), .C(n96), .D(\x[0][4] ), .Q(n279) );
  INV3 U366 ( .A(n278), .Q(n634) );
  AOI221 U367 ( .A(n115), .B(\x[1][5] ), .C(n96), .D(\x[0][5] ), .Q(n278) );
  INV3 U368 ( .A(n277), .Q(n635) );
  AOI221 U369 ( .A(n118), .B(\x[1][6] ), .C(n96), .D(\x[0][6] ), .Q(n277) );
  INV3 U370 ( .A(n276), .Q(n636) );
  AOI221 U371 ( .A(n120), .B(\x[1][7] ), .C(n96), .D(\x[0][7] ), .Q(n276) );
  INV3 U372 ( .A(n513), .Q(n125) );
  AOI221 U373 ( .A(n119), .B(\x[30][2] ), .C(n102), .D(\x[29][2] ), .Q(n513)
         );
  INV3 U374 ( .A(n497), .Q(n141) );
  AOI221 U375 ( .A(n117), .B(\x[28][2] ), .C(n110), .D(\x[27][2] ), .Q(n497)
         );
  INV3 U376 ( .A(n496), .Q(n142) );
  AOI221 U377 ( .A(n117), .B(\x[28][3] ), .C(n110), .D(\x[27][3] ), .Q(n496)
         );
  INV3 U378 ( .A(n495), .Q(n143) );
  AOI221 U379 ( .A(n117), .B(\x[28][4] ), .C(n110), .D(\x[27][4] ), .Q(n495)
         );
  INV3 U380 ( .A(n494), .Q(n144) );
  AOI221 U381 ( .A(n117), .B(\x[28][5] ), .C(n110), .D(\x[27][5] ), .Q(n494)
         );
  INV3 U382 ( .A(n493), .Q(n145) );
  AOI221 U383 ( .A(n117), .B(\x[28][6] ), .C(n110), .D(\x[27][6] ), .Q(n493)
         );
  INV3 U384 ( .A(n492), .Q(n146) );
  AOI221 U385 ( .A(n117), .B(\x[28][7] ), .C(n110), .D(\x[27][7] ), .Q(n492)
         );
  INV3 U386 ( .A(n491), .Q(n147) );
  AOI221 U387 ( .A(n117), .B(\x[27][0] ), .C(n110), .D(\x[26][0] ), .Q(n491)
         );
  INV3 U388 ( .A(n490), .Q(n148) );
  AOI221 U389 ( .A(n117), .B(\x[27][1] ), .C(n110), .D(\x[26][1] ), .Q(n490)
         );
  INV3 U390 ( .A(n489), .Q(n149) );
  AOI221 U391 ( .A(n117), .B(\x[27][2] ), .C(n109), .D(\x[26][2] ), .Q(n489)
         );
  INV3 U392 ( .A(n488), .Q(n150) );
  AOI221 U393 ( .A(n117), .B(\x[27][3] ), .C(n109), .D(\x[26][3] ), .Q(n488)
         );
  INV3 U394 ( .A(n487), .Q(n151) );
  AOI221 U395 ( .A(n117), .B(\x[27][4] ), .C(n109), .D(\x[26][4] ), .Q(n487)
         );
  INV3 U396 ( .A(n486), .Q(n152) );
  AOI221 U397 ( .A(n117), .B(\x[27][5] ), .C(n109), .D(\x[26][5] ), .Q(n486)
         );
  INV3 U398 ( .A(n485), .Q(n153) );
  AOI221 U399 ( .A(n117), .B(\x[27][6] ), .C(n109), .D(\x[26][6] ), .Q(n485)
         );
  INV3 U400 ( .A(n484), .Q(n154) );
  AOI221 U401 ( .A(n117), .B(\x[27][7] ), .C(n109), .D(\x[26][7] ), .Q(n484)
         );
  INV3 U402 ( .A(n483), .Q(n155) );
  AOI221 U403 ( .A(n117), .B(\x[26][0] ), .C(n109), .D(\x[25][0] ), .Q(n483)
         );
  INV3 U404 ( .A(n482), .Q(n156) );
  AOI221 U405 ( .A(n117), .B(\x[26][1] ), .C(n109), .D(\x[25][1] ), .Q(n482)
         );
  INV3 U406 ( .A(n481), .Q(n157) );
  AOI221 U407 ( .A(n117), .B(\x[26][2] ), .C(n109), .D(\x[25][2] ), .Q(n481)
         );
  INV3 U408 ( .A(n480), .Q(n158) );
  AOI221 U409 ( .A(n117), .B(\x[26][3] ), .C(n109), .D(\x[25][3] ), .Q(n480)
         );
  INV3 U410 ( .A(n479), .Q(n159) );
  AOI221 U411 ( .A(n117), .B(\x[26][4] ), .C(n109), .D(\x[25][4] ), .Q(n479)
         );
  INV3 U412 ( .A(n478), .Q(n160) );
  AOI221 U413 ( .A(n117), .B(\x[26][5] ), .C(n109), .D(\x[25][5] ), .Q(n478)
         );
  INV3 U414 ( .A(n477), .Q(n161) );
  AOI221 U415 ( .A(n117), .B(\x[26][6] ), .C(n109), .D(\x[25][6] ), .Q(n477)
         );
  INV3 U416 ( .A(n476), .Q(n162) );
  AOI221 U417 ( .A(n117), .B(\x[26][7] ), .C(n109), .D(\x[25][7] ), .Q(n476)
         );
  INV3 U418 ( .A(n453), .Q(n185) );
  AOI221 U419 ( .A(n119), .B(\x[23][6] ), .C(n107), .D(\x[22][6] ), .Q(n453)
         );
  INV3 U420 ( .A(n452), .Q(n186) );
  AOI221 U421 ( .A(n119), .B(\x[23][7] ), .C(n107), .D(\x[22][7] ), .Q(n452)
         );
  INV3 U422 ( .A(n451), .Q(n187) );
  AOI221 U423 ( .A(n119), .B(\x[22][0] ), .C(n107), .D(\x[21][0] ), .Q(n451)
         );
  INV3 U424 ( .A(n450), .Q(n188) );
  AOI221 U425 ( .A(n119), .B(\x[22][1] ), .C(n107), .D(\x[21][1] ), .Q(n450)
         );
  INV3 U426 ( .A(n449), .Q(n189) );
  AOI221 U427 ( .A(n119), .B(\x[22][2] ), .C(n107), .D(\x[21][2] ), .Q(n449)
         );
  INV3 U428 ( .A(n448), .Q(n190) );
  AOI221 U429 ( .A(n119), .B(\x[22][3] ), .C(n107), .D(\x[21][3] ), .Q(n448)
         );
  INV3 U430 ( .A(n447), .Q(n191) );
  AOI221 U431 ( .A(n119), .B(\x[22][4] ), .C(n107), .D(\x[21][4] ), .Q(n447)
         );
  INV3 U432 ( .A(n446), .Q(n192) );
  AOI221 U433 ( .A(n119), .B(\x[22][5] ), .C(n107), .D(\x[21][5] ), .Q(n446)
         );
  INV3 U434 ( .A(n445), .Q(n193) );
  AOI221 U435 ( .A(n119), .B(\x[22][6] ), .C(n107), .D(\x[21][6] ), .Q(n445)
         );
  INV3 U436 ( .A(n444), .Q(n194) );
  AOI221 U437 ( .A(n119), .B(\x[22][7] ), .C(n107), .D(\x[21][7] ), .Q(n444)
         );
  INV3 U438 ( .A(n443), .Q(n195) );
  AOI221 U439 ( .A(n119), .B(\x[21][0] ), .C(n107), .D(\x[20][0] ), .Q(n443)
         );
  INV3 U440 ( .A(n442), .Q(n196) );
  AOI221 U441 ( .A(n119), .B(\x[21][1] ), .C(n107), .D(\x[20][1] ), .Q(n442)
         );
  INV3 U442 ( .A(n441), .Q(n197) );
  AOI221 U443 ( .A(n119), .B(\x[21][2] ), .C(n106), .D(\x[20][2] ), .Q(n441)
         );
  INV3 U444 ( .A(n440), .Q(n198) );
  AOI221 U445 ( .A(n119), .B(\x[21][3] ), .C(n106), .D(\x[20][3] ), .Q(n440)
         );
  INV3 U446 ( .A(n439), .Q(n199) );
  AOI221 U447 ( .A(n119), .B(\x[21][4] ), .C(n106), .D(\x[20][4] ), .Q(n439)
         );
  INV3 U448 ( .A(n438), .Q(n200) );
  AOI221 U449 ( .A(n119), .B(\x[21][5] ), .C(n106), .D(\x[20][5] ), .Q(n438)
         );
  INV3 U450 ( .A(n437), .Q(n201) );
  AOI221 U451 ( .A(n119), .B(\x[21][6] ), .C(n106), .D(\x[20][6] ), .Q(n437)
         );
  INV3 U452 ( .A(n436), .Q(n202) );
  AOI221 U453 ( .A(n119), .B(\x[21][7] ), .C(n106), .D(\x[20][7] ), .Q(n436)
         );
  INV3 U454 ( .A(n435), .Q(n203) );
  AOI221 U455 ( .A(n119), .B(\x[20][0] ), .C(n106), .D(\x[19][0] ), .Q(n435)
         );
  INV3 U456 ( .A(n434), .Q(n204) );
  AOI221 U457 ( .A(n119), .B(\x[20][1] ), .C(n106), .D(\x[19][1] ), .Q(n434)
         );
  INV3 U458 ( .A(n433), .Q(n205) );
  AOI221 U459 ( .A(n119), .B(\x[20][2] ), .C(n106), .D(\x[19][2] ), .Q(n433)
         );
  INV3 U460 ( .A(n410), .Q(n228) );
  AOI221 U461 ( .A(n121), .B(\x[17][1] ), .C(n105), .D(\x[16][1] ), .Q(n410)
         );
  INV3 U462 ( .A(n409), .Q(n229) );
  AOI221 U463 ( .A(n121), .B(\x[17][2] ), .C(n104), .D(\x[16][2] ), .Q(n409)
         );
  INV3 U464 ( .A(n408), .Q(n230) );
  AOI221 U465 ( .A(n121), .B(\x[17][3] ), .C(n104), .D(\x[16][3] ), .Q(n408)
         );
  INV3 U466 ( .A(n407), .Q(n231) );
  AOI221 U467 ( .A(n121), .B(\x[17][4] ), .C(n104), .D(\x[16][4] ), .Q(n407)
         );
  INV3 U468 ( .A(n406), .Q(n232) );
  AOI221 U469 ( .A(n121), .B(\x[17][5] ), .C(n104), .D(\x[16][5] ), .Q(n406)
         );
  INV3 U470 ( .A(n405), .Q(n233) );
  AOI221 U471 ( .A(n121), .B(\x[17][6] ), .C(n104), .D(\x[16][6] ), .Q(n405)
         );
  INV3 U472 ( .A(n404), .Q(n234) );
  AOI221 U473 ( .A(n121), .B(\x[17][7] ), .C(n104), .D(\x[16][7] ), .Q(n404)
         );
  INV3 U474 ( .A(n403), .Q(n235) );
  AOI221 U475 ( .A(n121), .B(\x[16][0] ), .C(n104), .D(\x[15][0] ), .Q(n403)
         );
  INV3 U476 ( .A(n402), .Q(n236) );
  AOI221 U477 ( .A(n121), .B(\x[16][1] ), .C(n104), .D(\x[15][1] ), .Q(n402)
         );
  INV3 U478 ( .A(n401), .Q(n237) );
  AOI221 U479 ( .A(n121), .B(\x[16][2] ), .C(n104), .D(\x[15][2] ), .Q(n401)
         );
  INV3 U480 ( .A(n400), .Q(n238) );
  AOI221 U481 ( .A(n121), .B(\x[16][3] ), .C(n104), .D(\x[15][3] ), .Q(n400)
         );
  INV3 U482 ( .A(n399), .Q(n239) );
  AOI221 U483 ( .A(n121), .B(\x[16][4] ), .C(n104), .D(\x[15][4] ), .Q(n399)
         );
  INV3 U484 ( .A(n398), .Q(n240) );
  AOI221 U485 ( .A(n121), .B(\x[16][5] ), .C(n104), .D(\x[15][5] ), .Q(n398)
         );
  INV3 U486 ( .A(n397), .Q(n241) );
  AOI221 U487 ( .A(n121), .B(\x[16][6] ), .C(n104), .D(\x[15][6] ), .Q(n397)
         );
  INV3 U488 ( .A(n396), .Q(n242) );
  AOI221 U489 ( .A(n121), .B(\x[16][7] ), .C(n104), .D(\x[15][7] ), .Q(n396)
         );
  INV3 U490 ( .A(n395), .Q(n243) );
  AOI221 U491 ( .A(n121), .B(\x[15][0] ), .C(n104), .D(\x[14][0] ), .Q(n395)
         );
  INV3 U492 ( .A(n394), .Q(n244) );
  AOI221 U493 ( .A(n121), .B(\x[15][1] ), .C(n104), .D(\x[14][1] ), .Q(n394)
         );
  INV3 U494 ( .A(n393), .Q(n245) );
  AOI221 U495 ( .A(n121), .B(\x[15][2] ), .C(n103), .D(\x[14][2] ), .Q(n393)
         );
  INV3 U496 ( .A(n392), .Q(n246) );
  AOI221 U497 ( .A(n121), .B(\x[15][3] ), .C(n103), .D(\x[14][3] ), .Q(n392)
         );
  INV3 U498 ( .A(n391), .Q(n247) );
  AOI221 U499 ( .A(n121), .B(\x[15][4] ), .C(n103), .D(\x[14][4] ), .Q(n391)
         );
  INV3 U500 ( .A(n390), .Q(n248) );
  AOI221 U501 ( .A(n121), .B(\x[15][5] ), .C(n103), .D(\x[14][5] ), .Q(n390)
         );
  INV3 U502 ( .A(n389), .Q(n257) );
  AOI221 U503 ( .A(n121), .B(\x[15][6] ), .C(n103), .D(\x[14][6] ), .Q(n389)
         );
  INV3 U504 ( .A(n386), .Q(n526) );
  AOI221 U505 ( .A(n122), .B(\x[14][1] ), .C(n103), .D(\x[13][1] ), .Q(n386)
         );
  INV3 U506 ( .A(n349), .Q(n563) );
  AOI221 U507 ( .A(n95), .B(\x[10][6] ), .C(n101), .D(\x[9][6] ), .Q(n349) );
  INV3 U508 ( .A(n346), .Q(n566) );
  AOI221 U509 ( .A(n95), .B(\x[9][1] ), .C(n101), .D(\x[8][1] ), .Q(n346) );
  INV3 U510 ( .A(n345), .Q(n567) );
  AOI221 U511 ( .A(n259), .B(\x[9][2] ), .C(n100), .D(\x[8][2] ), .Q(n345) );
  INV3 U512 ( .A(n344), .Q(n568) );
  AOI221 U513 ( .A(n259), .B(\x[9][3] ), .C(n100), .D(\x[8][3] ), .Q(n344) );
  INV3 U514 ( .A(n343), .Q(n569) );
  AOI221 U515 ( .A(n259), .B(\x[9][4] ), .C(n100), .D(\x[8][4] ), .Q(n343) );
  INV3 U516 ( .A(n342), .Q(n570) );
  AOI221 U517 ( .A(n259), .B(\x[9][5] ), .C(n100), .D(\x[8][5] ), .Q(n342) );
  INV3 U518 ( .A(n341), .Q(n571) );
  AOI221 U519 ( .A(n259), .B(\x[9][6] ), .C(n100), .D(\x[8][6] ), .Q(n341) );
  INV3 U520 ( .A(n340), .Q(n572) );
  AOI221 U521 ( .A(n259), .B(\x[9][7] ), .C(n100), .D(\x[8][7] ), .Q(n340) );
  INV3 U522 ( .A(n339), .Q(n573) );
  AOI221 U523 ( .A(n259), .B(\x[8][0] ), .C(n100), .D(\x[7][0] ), .Q(n339) );
  INV3 U524 ( .A(n338), .Q(n574) );
  AOI221 U525 ( .A(n259), .B(\x[8][1] ), .C(n100), .D(\x[7][1] ), .Q(n338) );
  INV3 U526 ( .A(n337), .Q(n575) );
  AOI221 U527 ( .A(n259), .B(\x[8][2] ), .C(n100), .D(\x[7][2] ), .Q(n337) );
  INV3 U528 ( .A(n336), .Q(n576) );
  AOI221 U529 ( .A(n259), .B(\x[8][3] ), .C(n100), .D(\x[7][3] ), .Q(n336) );
  INV3 U530 ( .A(n335), .Q(n577) );
  AOI221 U531 ( .A(n259), .B(\x[8][4] ), .C(n100), .D(\x[7][4] ), .Q(n335) );
  INV3 U532 ( .A(n334), .Q(n578) );
  AOI221 U533 ( .A(n259), .B(\x[8][5] ), .C(n100), .D(\x[7][5] ), .Q(n334) );
  INV3 U534 ( .A(n333), .Q(n579) );
  AOI221 U535 ( .A(n259), .B(\x[8][6] ), .C(n100), .D(\x[7][6] ), .Q(n333) );
  INV3 U536 ( .A(n332), .Q(n580) );
  AOI221 U537 ( .A(n259), .B(\x[8][7] ), .C(n100), .D(\x[7][7] ), .Q(n332) );
  INV3 U538 ( .A(n331), .Q(n581) );
  AOI221 U539 ( .A(n259), .B(\x[7][0] ), .C(n100), .D(\x[6][0] ), .Q(n331) );
  INV3 U540 ( .A(n330), .Q(n582) );
  AOI221 U541 ( .A(n259), .B(\x[7][1] ), .C(n100), .D(\x[6][1] ), .Q(n330) );
  INV3 U542 ( .A(n329), .Q(n583) );
  AOI221 U543 ( .A(n259), .B(\x[7][2] ), .C(n99), .D(\x[6][2] ), .Q(n329) );
  INV3 U544 ( .A(n328), .Q(n584) );
  AOI221 U545 ( .A(n95), .B(\x[7][3] ), .C(n99), .D(\x[6][3] ), .Q(n328) );
  INV3 U546 ( .A(n327), .Q(n585) );
  AOI221 U547 ( .A(n95), .B(\x[7][4] ), .C(n99), .D(\x[6][4] ), .Q(n327) );
  INV3 U548 ( .A(n303), .Q(n609) );
  AOI221 U549 ( .A(n116), .B(\x[4][4] ), .C(n98), .D(\x[3][4] ), .Q(n303) );
  INV3 U550 ( .A(n302), .Q(n610) );
  AOI221 U551 ( .A(n116), .B(\x[4][5] ), .C(n98), .D(\x[3][5] ), .Q(n302) );
  INV3 U552 ( .A(n301), .Q(n611) );
  AOI221 U553 ( .A(n116), .B(\x[4][6] ), .C(n98), .D(\x[3][6] ), .Q(n301) );
  INV3 U554 ( .A(n300), .Q(n612) );
  AOI221 U555 ( .A(n116), .B(\x[4][7] ), .C(n98), .D(\x[3][7] ), .Q(n300) );
  INV3 U556 ( .A(n299), .Q(n613) );
  AOI221 U557 ( .A(n116), .B(\x[3][0] ), .C(n98), .D(\x[2][0] ), .Q(n299) );
  INV3 U558 ( .A(n298), .Q(n614) );
  AOI221 U559 ( .A(n116), .B(\x[3][1] ), .C(n98), .D(\x[2][1] ), .Q(n298) );
  INV3 U560 ( .A(n297), .Q(n615) );
  AOI221 U561 ( .A(n116), .B(\x[3][2] ), .C(n97), .D(\x[2][2] ), .Q(n297) );
  INV3 U562 ( .A(n296), .Q(n616) );
  AOI221 U563 ( .A(n116), .B(\x[3][3] ), .C(n97), .D(\x[2][3] ), .Q(n296) );
  INV3 U564 ( .A(n295), .Q(n617) );
  AOI221 U565 ( .A(n116), .B(\x[3][4] ), .C(n97), .D(\x[2][4] ), .Q(n295) );
  INV3 U566 ( .A(n294), .Q(n618) );
  AOI221 U567 ( .A(n116), .B(\x[3][5] ), .C(n97), .D(\x[2][5] ), .Q(n294) );
  INV3 U568 ( .A(n293), .Q(n619) );
  AOI221 U569 ( .A(n116), .B(\x[3][6] ), .C(n97), .D(\x[2][6] ), .Q(n293) );
  INV3 U570 ( .A(n292), .Q(n620) );
  AOI221 U571 ( .A(n116), .B(\x[3][7] ), .C(n97), .D(\x[2][7] ), .Q(n292) );
  INV3 U572 ( .A(n291), .Q(n621) );
  AOI221 U573 ( .A(n116), .B(\x[2][0] ), .C(n97), .D(\x[1][0] ), .Q(n291) );
  INV3 U574 ( .A(n290), .Q(n622) );
  AOI221 U575 ( .A(n116), .B(\x[2][1] ), .C(n97), .D(\x[1][1] ), .Q(n290) );
  INV3 U576 ( .A(n289), .Q(n623) );
  AOI221 U577 ( .A(n116), .B(\x[2][2] ), .C(n97), .D(\x[1][2] ), .Q(n289) );
  INV3 U578 ( .A(n288), .Q(n624) );
  AOI221 U579 ( .A(n116), .B(\x[2][3] ), .C(n97), .D(\x[1][3] ), .Q(n288) );
  INV3 U580 ( .A(n287), .Q(n625) );
  AOI221 U581 ( .A(n116), .B(\x[2][4] ), .C(n97), .D(\x[1][4] ), .Q(n287) );
  INV3 U582 ( .A(n286), .Q(n626) );
  AOI221 U583 ( .A(n116), .B(\x[2][5] ), .C(n97), .D(\x[1][5] ), .Q(n286) );
  INV3 U584 ( .A(n285), .Q(n627) );
  AOI221 U585 ( .A(n116), .B(\x[2][6] ), .C(n97), .D(\x[1][6] ), .Q(n285) );
  INV3 U586 ( .A(n284), .Q(n628) );
  AOI221 U587 ( .A(n116), .B(\x[2][7] ), .C(n97), .D(\x[1][7] ), .Q(n284) );
  INV3 U588 ( .A(n283), .Q(n629) );
  AOI221 U589 ( .A(n116), .B(\x[1][0] ), .C(n97), .D(\x[0][0] ), .Q(n283) );
  INV3 U590 ( .A(n282), .Q(n630) );
  AOI221 U591 ( .A(n116), .B(\x[1][1] ), .C(n97), .D(\x[0][1] ), .Q(n282) );
  INV3 U592 ( .A(n514), .Q(n124) );
  AOI221 U593 ( .A(n116), .B(\x[30][1] ), .C(n110), .D(\x[29][1] ), .Q(n514)
         );
  INV3 U594 ( .A(n385), .Q(n527) );
  AOI221 U595 ( .A(n122), .B(\x[14][2] ), .C(n103), .D(\x[13][2] ), .Q(n385)
         );
  INV3 U596 ( .A(n384), .Q(n528) );
  AOI221 U597 ( .A(n120), .B(\x[14][3] ), .C(n103), .D(\x[13][3] ), .Q(n384)
         );
  INV3 U598 ( .A(n383), .Q(n529) );
  AOI221 U599 ( .A(n122), .B(\x[14][4] ), .C(n103), .D(\x[13][4] ), .Q(n383)
         );
  INV3 U600 ( .A(n382), .Q(n530) );
  AOI221 U601 ( .A(n122), .B(\x[14][5] ), .C(n103), .D(\x[13][5] ), .Q(n382)
         );
  INV3 U602 ( .A(n381), .Q(n531) );
  AOI221 U603 ( .A(n122), .B(\x[14][6] ), .C(n103), .D(\x[13][6] ), .Q(n381)
         );
  INV3 U604 ( .A(n380), .Q(n532) );
  AOI221 U605 ( .A(n122), .B(\x[14][7] ), .C(n103), .D(\x[13][7] ), .Q(n380)
         );
  INV3 U606 ( .A(n379), .Q(n533) );
  AOI221 U607 ( .A(n122), .B(\x[13][0] ), .C(n103), .D(\x[12][0] ), .Q(n379)
         );
  INV3 U608 ( .A(n378), .Q(n534) );
  AOI221 U609 ( .A(n122), .B(\x[13][1] ), .C(n103), .D(\x[12][1] ), .Q(n378)
         );
  INV3 U610 ( .A(n377), .Q(n535) );
  AOI221 U611 ( .A(n122), .B(\x[13][2] ), .C(n102), .D(\x[12][2] ), .Q(n377)
         );
  INV3 U612 ( .A(n376), .Q(n536) );
  AOI221 U613 ( .A(n122), .B(\x[13][3] ), .C(n102), .D(\x[12][3] ), .Q(n376)
         );
  INV3 U614 ( .A(n375), .Q(n537) );
  AOI221 U615 ( .A(n122), .B(\x[13][4] ), .C(n102), .D(\x[12][4] ), .Q(n375)
         );
  INV3 U616 ( .A(n374), .Q(n538) );
  AOI221 U617 ( .A(n122), .B(\x[13][5] ), .C(n102), .D(\x[12][5] ), .Q(n374)
         );
  INV3 U618 ( .A(n372), .Q(n540) );
  AOI221 U619 ( .A(n122), .B(\x[13][7] ), .C(n102), .D(\x[12][7] ), .Q(n372)
         );
  INV3 U620 ( .A(n371), .Q(n541) );
  AOI221 U621 ( .A(n122), .B(\x[12][0] ), .C(n102), .D(\x[11][0] ), .Q(n371)
         );
  INV3 U622 ( .A(n370), .Q(n542) );
  AOI221 U623 ( .A(n122), .B(\x[12][1] ), .C(n102), .D(\x[11][1] ), .Q(n370)
         );
  INV3 U624 ( .A(n369), .Q(n543) );
  AOI221 U625 ( .A(n122), .B(\x[12][2] ), .C(n102), .D(\x[11][2] ), .Q(n369)
         );
  INV3 U626 ( .A(n515), .Q(n123) );
  AOI221 U627 ( .A(\x[30][0] ), .B(n114), .C(n109), .D(\x[29][0] ), .Q(n515)
         );
  INV3 U628 ( .A(n275), .Q(n637) );
  AOI221 U629 ( .A(Delay_Line_in[0]), .B(n96), .C(\x[0][0] ), .D(n117), .Q(
        n275) );
  INV3 U630 ( .A(n274), .Q(n638) );
  AOI221 U631 ( .A(Delay_Line_in[1]), .B(n96), .C(\x[0][1] ), .D(n114), .Q(
        n274) );
  INV3 U632 ( .A(n273), .Q(n639) );
  AOI221 U633 ( .A(Delay_Line_in[2]), .B(n96), .C(\x[0][2] ), .D(n119), .Q(
        n273) );
  INV3 U634 ( .A(n272), .Q(n640) );
  AOI221 U635 ( .A(Delay_Line_in[3]), .B(n96), .C(\x[0][3] ), .D(n121), .Q(
        n272) );
  INV3 U636 ( .A(n271), .Q(n641) );
  AOI221 U637 ( .A(Delay_Line_in[4]), .B(n96), .C(\x[0][4] ), .D(n114), .Q(
        n271) );
  INV3 U638 ( .A(n270), .Q(n642) );
  AOI221 U639 ( .A(Delay_Line_in[5]), .B(n96), .C(\x[0][5] ), .D(n116), .Q(
        n270) );
  INV3 U640 ( .A(n269), .Q(n643) );
  AOI221 U641 ( .A(Delay_Line_in[6]), .B(n96), .C(\x[0][6] ), .D(n114), .Q(
        n269) );
  INV3 U642 ( .A(n268), .Q(n644) );
  AOI221 U643 ( .A(Delay_Line_in[7]), .B(n96), .C(\x[0][7] ), .D(n114), .Q(
        n268) );
  NAND22 U644 ( .A(\x[31][0] ), .B(n114), .Q(n258) );
  NAND22 U645 ( .A(\x[31][1] ), .B(n114), .Q(n260) );
  NAND22 U646 ( .A(\x[31][2] ), .B(n114), .Q(n261) );
endmodule


module coeff_ram ( CLK, RESET, data_in, data_out, address, wb );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] address;
  input CLK, RESET, wb;
  wire   N10, N11, N12, N13, N14, \ram[0][7] , \ram[0][6] , \ram[0][5] ,
         \ram[0][4] , \ram[0][3] , \ram[0][2] , \ram[0][1] , \ram[0][0] ,
         \ram[1][7] , \ram[1][6] , \ram[1][5] , \ram[1][4] , \ram[1][3] ,
         \ram[1][2] , \ram[1][1] , \ram[1][0] , \ram[2][7] , \ram[2][6] ,
         \ram[2][5] , \ram[2][4] , \ram[2][3] , \ram[2][2] , \ram[2][1] ,
         \ram[2][0] , \ram[3][7] , \ram[3][6] , \ram[3][5] , \ram[3][4] ,
         \ram[3][3] , \ram[3][2] , \ram[3][1] , \ram[3][0] , \ram[4][7] ,
         \ram[4][6] , \ram[4][5] , \ram[4][4] , \ram[4][3] , \ram[4][2] ,
         \ram[4][1] , \ram[4][0] , \ram[5][7] , \ram[5][6] , \ram[5][5] ,
         \ram[5][4] , \ram[5][3] , \ram[5][2] , \ram[5][1] , \ram[5][0] ,
         \ram[6][7] , \ram[6][6] , \ram[6][5] , \ram[6][4] , \ram[6][3] ,
         \ram[6][2] , \ram[6][1] , \ram[6][0] , \ram[7][7] , \ram[7][6] ,
         \ram[7][5] , \ram[7][4] , \ram[7][3] , \ram[7][2] , \ram[7][1] ,
         \ram[7][0] , \ram[8][7] , \ram[8][6] , \ram[8][5] , \ram[8][4] ,
         \ram[8][3] , \ram[8][2] , \ram[8][1] , \ram[8][0] , \ram[9][7] ,
         \ram[9][6] , \ram[9][5] , \ram[9][4] , \ram[9][3] , \ram[9][2] ,
         \ram[9][1] , \ram[9][0] , \ram[10][7] , \ram[10][6] , \ram[10][5] ,
         \ram[10][4] , \ram[10][3] , \ram[10][2] , \ram[10][1] , \ram[10][0] ,
         \ram[11][7] , \ram[11][6] , \ram[11][5] , \ram[11][4] , \ram[11][3] ,
         \ram[11][2] , \ram[11][1] , \ram[11][0] , \ram[12][7] , \ram[12][6] ,
         \ram[12][5] , \ram[12][4] , \ram[12][3] , \ram[12][2] , \ram[12][1] ,
         \ram[12][0] , \ram[13][7] , \ram[13][6] , \ram[13][5] , \ram[13][4] ,
         \ram[13][3] , \ram[13][2] , \ram[13][1] , \ram[13][0] , \ram[14][7] ,
         \ram[14][6] , \ram[14][5] , \ram[14][4] , \ram[14][3] , \ram[14][2] ,
         \ram[14][1] , \ram[14][0] , \ram[15][7] , \ram[15][6] , \ram[15][5] ,
         \ram[15][4] , \ram[15][3] , \ram[15][2] , \ram[15][1] , \ram[15][0] ,
         \ram[16][7] , \ram[16][6] , \ram[16][5] , \ram[16][4] , \ram[16][3] ,
         \ram[16][2] , \ram[16][1] , \ram[16][0] , \ram[17][7] , \ram[17][6] ,
         \ram[17][5] , \ram[17][4] , \ram[17][3] , \ram[17][2] , \ram[17][1] ,
         \ram[17][0] , \ram[18][7] , \ram[18][6] , \ram[18][5] , \ram[18][4] ,
         \ram[18][3] , \ram[18][2] , \ram[18][1] , \ram[18][0] , \ram[19][7] ,
         \ram[19][6] , \ram[19][5] , \ram[19][4] , \ram[19][3] , \ram[19][2] ,
         \ram[19][1] , \ram[19][0] , \ram[20][7] , \ram[20][6] , \ram[20][5] ,
         \ram[20][4] , \ram[20][3] , \ram[20][2] , \ram[20][1] , \ram[20][0] ,
         \ram[21][7] , \ram[21][6] , \ram[21][5] , \ram[21][4] , \ram[21][3] ,
         \ram[21][2] , \ram[21][1] , \ram[21][0] , \ram[22][7] , \ram[22][6] ,
         \ram[22][5] , \ram[22][4] , \ram[22][3] , \ram[22][2] , \ram[22][1] ,
         \ram[22][0] , \ram[23][7] , \ram[23][6] , \ram[23][5] , \ram[23][4] ,
         \ram[23][3] , \ram[23][2] , \ram[23][1] , \ram[23][0] , \ram[24][7] ,
         \ram[24][6] , \ram[24][5] , \ram[24][4] , \ram[24][3] , \ram[24][2] ,
         \ram[24][1] , \ram[24][0] , \ram[25][7] , \ram[25][6] , \ram[25][5] ,
         \ram[25][4] , \ram[25][3] , \ram[25][2] , \ram[25][1] , \ram[25][0] ,
         \ram[26][7] , \ram[26][6] , \ram[26][5] , \ram[26][4] , \ram[26][3] ,
         \ram[26][2] , \ram[26][1] , \ram[26][0] , \ram[27][7] , \ram[27][6] ,
         \ram[27][5] , \ram[27][4] , \ram[27][3] , \ram[27][2] , \ram[27][1] ,
         \ram[27][0] , \ram[28][7] , \ram[28][6] , \ram[28][5] , \ram[28][4] ,
         \ram[28][3] , \ram[28][2] , \ram[28][1] , \ram[28][0] , \ram[29][7] ,
         \ram[29][6] , \ram[29][5] , \ram[29][4] , \ram[29][3] , \ram[29][2] ,
         \ram[29][1] , \ram[29][0] , \ram[30][7] , \ram[30][6] , \ram[30][5] ,
         \ram[30][4] , \ram[30][3] , \ram[30][2] , \ram[30][1] , \ram[30][0] ,
         \ram[31][7] , \ram[31][6] , \ram[31][5] , \ram[31][4] , \ram[31][3] ,
         \ram[31][2] , \ram[31][1] , \ram[31][0] , n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251;
  assign N10 = address[0];
  assign N11 = address[1];
  assign N12 = address[2];
  assign N13 = address[3];
  assign N14 = address[4];

  DFEC1 \ram_reg[2][7]  ( .D(n216), .E(n237), .C(CLK), .RN(n165), .Q(
        \ram[2][7] ) );
  DFEC1 \ram_reg[2][6]  ( .D(n212), .E(n237), .C(CLK), .RN(n165), .Q(
        \ram[2][6] ) );
  DFEC1 \ram_reg[6][7]  ( .D(n216), .E(n245), .C(CLK), .RN(n167), .Q(
        \ram[6][7] ) );
  DFEC1 \ram_reg[6][6]  ( .D(n212), .E(n245), .C(CLK), .RN(n167), .Q(
        \ram[6][6] ) );
  DFEC1 \ram_reg[10][7]  ( .D(n215), .E(n238), .C(CLK), .RN(n169), .Q(
        \ram[10][7] ) );
  DFEC1 \ram_reg[10][6]  ( .D(n211), .E(n238), .C(CLK), .RN(n169), .Q(
        \ram[10][6] ) );
  DFEC1 \ram_reg[14][7]  ( .D(n215), .E(n246), .C(CLK), .RN(n163), .Q(
        \ram[14][7] ) );
  DFEC1 \ram_reg[14][6]  ( .D(n211), .E(n246), .C(CLK), .RN(n162), .Q(
        \ram[14][6] ) );
  DFEC1 \ram_reg[22][7]  ( .D(n214), .E(n247), .C(CLK), .RN(n159), .Q(
        \ram[22][7] ) );
  DFEC1 \ram_reg[22][6]  ( .D(n210), .E(n247), .C(CLK), .RN(n159), .Q(
        \ram[22][6] ) );
  DFEC1 \ram_reg[26][7]  ( .D(n213), .E(n240), .C(CLK), .RN(n157), .Q(
        \ram[26][7] ) );
  DFEC1 \ram_reg[26][6]  ( .D(n209), .E(n240), .C(CLK), .RN(n157), .Q(
        \ram[26][6] ) );
  DFEC1 \ram_reg[30][7]  ( .D(n213), .E(n248), .C(CLK), .RN(n155), .Q(
        \ram[30][7] ) );
  DFEC1 \ram_reg[30][6]  ( .D(n209), .E(n248), .C(CLK), .RN(n155), .Q(
        \ram[30][6] ) );
  DFEP1 \ram_reg[18][7]  ( .D(n214), .E(n239), .C(CLK), .SN(n180), .Q(
        \ram[18][7] ) );
  DFEP1 \ram_reg[18][6]  ( .D(n210), .E(n239), .C(CLK), .SN(n180), .Q(
        \ram[18][6] ) );
  DFEC1 \ram_reg[0][7]  ( .D(n216), .E(n233), .C(CLK), .RN(n154), .Q(
        \ram[0][7] ) );
  DFEC1 \ram_reg[0][6]  ( .D(n212), .E(n233), .C(CLK), .RN(n166), .Q(
        \ram[0][6] ) );
  DFEC1 \ram_reg[1][7]  ( .D(n216), .E(n229), .C(CLK), .RN(n164), .Q(
        \ram[1][7] ) );
  DFEC1 \ram_reg[1][6]  ( .D(n212), .E(n229), .C(CLK), .RN(n165), .Q(
        \ram[1][6] ) );
  DFEC1 \ram_reg[5][7]  ( .D(n216), .E(n221), .C(CLK), .RN(n166), .Q(
        \ram[5][7] ) );
  DFEC1 \ram_reg[5][6]  ( .D(n212), .E(n221), .C(CLK), .RN(n166), .Q(
        \ram[5][6] ) );
  DFEC1 \ram_reg[9][7]  ( .D(n215), .E(n230), .C(CLK), .RN(n168), .Q(
        \ram[9][7] ) );
  DFEC1 \ram_reg[9][6]  ( .D(n211), .E(n230), .C(CLK), .RN(n169), .Q(
        \ram[9][6] ) );
  DFEC1 \ram_reg[11][7]  ( .D(n215), .E(n226), .C(CLK), .RN(n169), .Q(
        \ram[11][7] ) );
  DFEC1 \ram_reg[11][6]  ( .D(n211), .E(n226), .C(CLK), .RN(n169), .Q(
        \ram[11][6] ) );
  DFEC1 \ram_reg[15][7]  ( .D(n215), .E(n218), .C(CLK), .RN(n162), .Q(
        \ram[15][7] ) );
  DFEC1 \ram_reg[16][7]  ( .D(n214), .E(n235), .C(CLK), .RN(n162), .Q(
        \ram[16][7] ) );
  DFEC1 \ram_reg[17][7]  ( .D(n214), .E(n231), .C(CLK), .RN(n161), .Q(
        \ram[17][7] ) );
  DFEC1 \ram_reg[17][6]  ( .D(n210), .E(n231), .C(CLK), .RN(n161), .Q(
        \ram[17][6] ) );
  DFEC1 \ram_reg[20][7]  ( .D(n214), .E(n243), .C(CLK), .RN(n160), .Q(
        \ram[20][7] ) );
  DFEC1 \ram_reg[20][6]  ( .D(n210), .E(n243), .C(CLK), .RN(n160), .Q(
        \ram[20][6] ) );
  DFEC1 \ram_reg[21][7]  ( .D(n214), .E(n223), .C(CLK), .RN(n159), .Q(
        \ram[21][7] ) );
  DFEC1 \ram_reg[21][6]  ( .D(n210), .E(n223), .C(CLK), .RN(n159), .Q(
        \ram[21][6] ) );
  DFEC1 \ram_reg[25][7]  ( .D(n213), .E(n232), .C(CLK), .RN(n158), .Q(
        \ram[25][7] ) );
  DFEC1 \ram_reg[25][6]  ( .D(n209), .E(n232), .C(CLK), .RN(n157), .Q(
        \ram[25][6] ) );
  DFEC1 \ram_reg[29][7]  ( .D(n213), .E(n224), .C(CLK), .RN(n156), .Q(
        \ram[29][7] ) );
  DFEC1 \ram_reg[29][6]  ( .D(n209), .E(n224), .C(CLK), .RN(n156), .Q(
        \ram[29][6] ) );
  DFEC1 \ram_reg[31][7]  ( .D(n213), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][7] ) );
  DFEC1 \ram_reg[31][6]  ( .D(n209), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][6] ) );
  DFEP1 \ram_reg[3][7]  ( .D(n216), .E(n225), .C(CLK), .SN(n173), .Q(
        \ram[3][7] ) );
  DFEP1 \ram_reg[3][6]  ( .D(n212), .E(n225), .C(CLK), .SN(n173), .Q(
        \ram[3][6] ) );
  DFEP1 \ram_reg[4][7]  ( .D(n216), .E(n241), .C(CLK), .SN(n174), .Q(
        \ram[4][7] ) );
  DFEP1 \ram_reg[4][6]  ( .D(n212), .E(n241), .C(CLK), .SN(n174), .Q(
        \ram[4][6] ) );
  DFEP1 \ram_reg[7][7]  ( .D(n216), .E(n217), .C(CLK), .SN(n178), .Q(
        \ram[7][7] ) );
  DFEP1 \ram_reg[7][6]  ( .D(n212), .E(n217), .C(CLK), .SN(n178), .Q(
        \ram[7][6] ) );
  DFEP1 \ram_reg[8][7]  ( .D(n215), .E(n234), .C(CLK), .SN(n179), .Q(
        \ram[8][7] ) );
  DFEP1 \ram_reg[8][6]  ( .D(n211), .E(n234), .C(CLK), .SN(n179), .Q(
        \ram[8][6] ) );
  DFEP1 \ram_reg[12][7]  ( .D(n215), .E(n242), .C(CLK), .SN(n171), .Q(
        \ram[12][7] ) );
  DFEP1 \ram_reg[12][6]  ( .D(n211), .E(n242), .C(CLK), .SN(n170), .Q(
        \ram[12][6] ) );
  DFEP1 \ram_reg[13][7]  ( .D(n215), .E(n222), .C(CLK), .SN(n171), .Q(
        \ram[13][7] ) );
  DFEP1 \ram_reg[13][6]  ( .D(n211), .E(n222), .C(CLK), .SN(n171), .Q(
        \ram[13][6] ) );
  DFEP1 \ram_reg[15][6]  ( .D(n211), .E(n218), .C(CLK), .SN(n177), .Q(
        \ram[15][6] ) );
  DFEP1 \ram_reg[16][6]  ( .D(n210), .E(n235), .C(CLK), .SN(n179), .Q(
        \ram[16][6] ) );
  DFEP1 \ram_reg[19][7]  ( .D(n214), .E(n227), .C(CLK), .SN(n179), .Q(
        \ram[19][7] ) );
  DFEP1 \ram_reg[19][6]  ( .D(n210), .E(n227), .C(CLK), .SN(n179), .Q(
        \ram[19][6] ) );
  DFEP1 \ram_reg[23][7]  ( .D(n214), .E(n219), .C(CLK), .SN(n176), .Q(
        \ram[23][7] ) );
  DFEP1 \ram_reg[23][6]  ( .D(n210), .E(n219), .C(CLK), .SN(n176), .Q(
        \ram[23][6] ) );
  DFEP1 \ram_reg[24][7]  ( .D(n213), .E(n236), .C(CLK), .SN(n176), .Q(
        \ram[24][7] ) );
  DFEP1 \ram_reg[24][6]  ( .D(n209), .E(n236), .C(CLK), .SN(n175), .Q(
        \ram[24][6] ) );
  DFEP1 \ram_reg[27][7]  ( .D(n213), .E(n228), .C(CLK), .SN(n173), .Q(
        \ram[27][7] ) );
  DFEP1 \ram_reg[27][6]  ( .D(n209), .E(n228), .C(CLK), .SN(n173), .Q(
        \ram[27][6] ) );
  DFEP1 \ram_reg[28][7]  ( .D(n213), .E(n244), .C(CLK), .SN(n172), .Q(
        \ram[28][7] ) );
  DFEP1 \ram_reg[28][6]  ( .D(n209), .E(n244), .C(CLK), .SN(n175), .Q(
        \ram[28][6] ) );
  DFEC1 \ram_reg[2][5]  ( .D(n208), .E(n237), .C(CLK), .RN(n165), .Q(
        \ram[2][5] ) );
  DFEC1 \ram_reg[2][4]  ( .D(n204), .E(n237), .C(CLK), .RN(n168), .Q(
        \ram[2][4] ) );
  DFEC1 \ram_reg[6][5]  ( .D(n208), .E(n245), .C(CLK), .RN(n167), .Q(
        \ram[6][5] ) );
  DFEC1 \ram_reg[6][4]  ( .D(n204), .E(n245), .C(CLK), .RN(n167), .Q(
        \ram[6][4] ) );
  DFEC1 \ram_reg[10][5]  ( .D(n207), .E(n238), .C(CLK), .RN(n169), .Q(
        \ram[10][5] ) );
  DFEC1 \ram_reg[10][4]  ( .D(n203), .E(n238), .C(CLK), .RN(n169), .Q(
        \ram[10][4] ) );
  DFEC1 \ram_reg[14][4]  ( .D(n203), .E(n246), .C(CLK), .RN(n162), .Q(
        \ram[14][4] ) );
  DFEC1 \ram_reg[22][5]  ( .D(n206), .E(n247), .C(CLK), .RN(n159), .Q(
        \ram[22][5] ) );
  DFEC1 \ram_reg[22][4]  ( .D(n202), .E(n247), .C(CLK), .RN(n158), .Q(
        \ram[22][4] ) );
  DFEC1 \ram_reg[26][5]  ( .D(n205), .E(n240), .C(CLK), .RN(n157), .Q(
        \ram[26][5] ) );
  DFEC1 \ram_reg[26][4]  ( .D(n201), .E(n240), .C(CLK), .RN(n157), .Q(
        \ram[26][4] ) );
  DFEC1 \ram_reg[30][5]  ( .D(n205), .E(n248), .C(CLK), .RN(n155), .Q(
        \ram[30][5] ) );
  DFEC1 \ram_reg[30][4]  ( .D(n201), .E(n248), .C(CLK), .RN(n155), .Q(
        \ram[30][4] ) );
  DFEP1 \ram_reg[14][5]  ( .D(n207), .E(n246), .C(CLK), .SN(n175), .Q(
        \ram[14][5] ) );
  DFEP1 \ram_reg[18][5]  ( .D(n206), .E(n239), .C(CLK), .SN(n180), .Q(
        \ram[18][5] ) );
  DFEP1 \ram_reg[18][4]  ( .D(n202), .E(n239), .C(CLK), .SN(n180), .Q(
        \ram[18][4] ) );
  DFEC1 \ram_reg[0][5]  ( .D(n208), .E(n233), .C(CLK), .RN(n164), .Q(
        \ram[0][5] ) );
  DFEC1 \ram_reg[0][4]  ( .D(n204), .E(n233), .C(CLK), .RN(n164), .Q(
        \ram[0][4] ) );
  DFEC1 \ram_reg[1][5]  ( .D(n208), .E(n229), .C(CLK), .RN(n165), .Q(
        \ram[1][5] ) );
  DFEC1 \ram_reg[1][4]  ( .D(n204), .E(n229), .C(CLK), .RN(n165), .Q(
        \ram[1][4] ) );
  DFEC1 \ram_reg[5][5]  ( .D(n208), .E(n221), .C(CLK), .RN(n166), .Q(
        \ram[5][5] ) );
  DFEC1 \ram_reg[5][4]  ( .D(n204), .E(n221), .C(CLK), .RN(n167), .Q(
        \ram[5][4] ) );
  DFEC1 \ram_reg[9][5]  ( .D(n207), .E(n230), .C(CLK), .RN(n170), .Q(
        \ram[9][5] ) );
  DFEC1 \ram_reg[9][4]  ( .D(n203), .E(n230), .C(CLK), .RN(n170), .Q(
        \ram[9][4] ) );
  DFEC1 \ram_reg[11][5]  ( .D(n207), .E(n226), .C(CLK), .RN(n168), .Q(
        \ram[11][5] ) );
  DFEC1 \ram_reg[11][4]  ( .D(n203), .E(n226), .C(CLK), .RN(n169), .Q(
        \ram[11][4] ) );
  DFEC1 \ram_reg[12][4]  ( .D(n203), .E(n242), .C(CLK), .RN(n163), .Q(
        \ram[12][4] ) );
  DFEC1 \ram_reg[15][4]  ( .D(n203), .E(n218), .C(CLK), .RN(n162), .Q(
        \ram[15][4] ) );
  DFEC1 \ram_reg[16][4]  ( .D(n202), .E(n235), .C(CLK), .RN(n162), .Q(
        \ram[16][4] ) );
  DFEC1 \ram_reg[17][4]  ( .D(n202), .E(n231), .C(CLK), .RN(n161), .Q(
        \ram[17][4] ) );
  DFEC1 \ram_reg[19][4]  ( .D(n202), .E(n227), .C(CLK), .RN(n160), .Q(
        \ram[19][4] ) );
  DFEC1 \ram_reg[20][5]  ( .D(n206), .E(n243), .C(CLK), .RN(n160), .Q(
        \ram[20][5] ) );
  DFEC1 \ram_reg[20][4]  ( .D(n202), .E(n243), .C(CLK), .RN(n160), .Q(
        \ram[20][4] ) );
  DFEC1 \ram_reg[21][5]  ( .D(n206), .E(n223), .C(CLK), .RN(n159), .Q(
        \ram[21][5] ) );
  DFEC1 \ram_reg[21][4]  ( .D(n202), .E(n223), .C(CLK), .RN(n159), .Q(
        \ram[21][4] ) );
  DFEC1 \ram_reg[25][5]  ( .D(n205), .E(n232), .C(CLK), .RN(n157), .Q(
        \ram[25][5] ) );
  DFEC1 \ram_reg[25][4]  ( .D(n201), .E(n232), .C(CLK), .RN(n157), .Q(
        \ram[25][4] ) );
  DFEC1 \ram_reg[29][5]  ( .D(n205), .E(n224), .C(CLK), .RN(n156), .Q(
        \ram[29][5] ) );
  DFEC1 \ram_reg[29][4]  ( .D(n201), .E(n224), .C(CLK), .RN(n156), .Q(
        \ram[29][4] ) );
  DFEC1 \ram_reg[31][5]  ( .D(n205), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][5] ) );
  DFEC1 \ram_reg[31][4]  ( .D(n201), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][4] ) );
  DFEP1 \ram_reg[3][5]  ( .D(n208), .E(n225), .C(CLK), .SN(n173), .Q(
        \ram[3][5] ) );
  DFEP1 \ram_reg[3][4]  ( .D(n204), .E(n225), .C(CLK), .SN(n173), .Q(
        \ram[3][4] ) );
  DFEP1 \ram_reg[4][5]  ( .D(n208), .E(n241), .C(CLK), .SN(n174), .Q(
        \ram[4][5] ) );
  DFEP1 \ram_reg[4][4]  ( .D(n204), .E(n241), .C(CLK), .SN(n174), .Q(
        \ram[4][4] ) );
  DFEP1 \ram_reg[7][5]  ( .D(n208), .E(n217), .C(CLK), .SN(n178), .Q(
        \ram[7][5] ) );
  DFEP1 \ram_reg[7][4]  ( .D(n204), .E(n217), .C(CLK), .SN(n178), .Q(
        \ram[7][4] ) );
  DFEP1 \ram_reg[8][5]  ( .D(n207), .E(n234), .C(CLK), .SN(n179), .Q(
        \ram[8][5] ) );
  DFEP1 \ram_reg[8][4]  ( .D(n203), .E(n234), .C(CLK), .SN(n180), .Q(
        \ram[8][4] ) );
  DFEP1 \ram_reg[12][5]  ( .D(n207), .E(n242), .C(CLK), .SN(n171), .Q(
        \ram[12][5] ) );
  DFEP1 \ram_reg[13][5]  ( .D(n207), .E(n222), .C(CLK), .SN(n172), .Q(
        \ram[13][5] ) );
  DFEP1 \ram_reg[13][4]  ( .D(n203), .E(n222), .C(CLK), .SN(n172), .Q(
        \ram[13][4] ) );
  DFEP1 \ram_reg[15][5]  ( .D(n207), .E(n218), .C(CLK), .SN(n177), .Q(
        \ram[15][5] ) );
  DFEP1 \ram_reg[16][5]  ( .D(n206), .E(n235), .C(CLK), .SN(n181), .Q(
        \ram[16][5] ) );
  DFEP1 \ram_reg[17][5]  ( .D(n206), .E(n231), .C(CLK), .SN(n180), .Q(
        \ram[17][5] ) );
  DFEP1 \ram_reg[19][5]  ( .D(n206), .E(n227), .C(CLK), .SN(n179), .Q(
        \ram[19][5] ) );
  DFEP1 \ram_reg[23][5]  ( .D(n206), .E(n219), .C(CLK), .SN(n176), .Q(
        \ram[23][5] ) );
  DFEP1 \ram_reg[23][4]  ( .D(n202), .E(n219), .C(CLK), .SN(n176), .Q(
        \ram[23][4] ) );
  DFEP1 \ram_reg[24][5]  ( .D(n205), .E(n236), .C(CLK), .SN(n175), .Q(
        \ram[24][5] ) );
  DFEP1 \ram_reg[24][4]  ( .D(n201), .E(n236), .C(CLK), .SN(n175), .Q(
        \ram[24][4] ) );
  DFEP1 \ram_reg[27][5]  ( .D(n205), .E(n228), .C(CLK), .SN(n173), .Q(
        \ram[27][5] ) );
  DFEP1 \ram_reg[27][4]  ( .D(n201), .E(n228), .C(CLK), .SN(n173), .Q(
        \ram[27][4] ) );
  DFEP1 \ram_reg[28][5]  ( .D(n205), .E(n244), .C(CLK), .SN(n172), .Q(
        \ram[28][5] ) );
  DFEP1 \ram_reg[28][4]  ( .D(n201), .E(n244), .C(CLK), .SN(n172), .Q(
        \ram[28][4] ) );
  DFEC1 \ram_reg[2][3]  ( .D(n200), .E(n237), .C(CLK), .RN(n166), .Q(
        \ram[2][3] ) );
  DFEC1 \ram_reg[6][3]  ( .D(n200), .E(n245), .C(CLK), .RN(n167), .Q(
        \ram[6][3] ) );
  DFEC1 \ram_reg[18][3]  ( .D(n198), .E(n239), .C(CLK), .RN(n161), .Q(
        \ram[18][3] ) );
  DFEC1 \ram_reg[22][3]  ( .D(n198), .E(n247), .C(CLK), .RN(n158), .Q(
        \ram[22][3] ) );
  DFEC1 \ram_reg[26][3]  ( .D(n197), .E(n240), .C(CLK), .RN(n156), .Q(
        \ram[26][3] ) );
  DFEC1 \ram_reg[30][3]  ( .D(n197), .E(n248), .C(CLK), .RN(n155), .Q(
        \ram[30][3] ) );
  DFEP1 \ram_reg[10][3]  ( .D(n199), .E(n238), .C(CLK), .SN(n171), .Q(
        \ram[10][3] ) );
  DFEP1 \ram_reg[14][3]  ( .D(n199), .E(n246), .C(CLK), .SN(n176), .Q(
        \ram[14][3] ) );
  DFEC1 \ram_reg[0][3]  ( .D(n200), .E(n233), .C(CLK), .RN(n164), .Q(
        \ram[0][3] ) );
  DFEC1 \ram_reg[1][3]  ( .D(n200), .E(n229), .C(CLK), .RN(n165), .Q(
        \ram[1][3] ) );
  DFEC1 \ram_reg[5][3]  ( .D(n200), .E(n221), .C(CLK), .RN(n167), .Q(
        \ram[5][3] ) );
  DFEC1 \ram_reg[9][3]  ( .D(n199), .E(n230), .C(CLK), .RN(n170), .Q(
        \ram[9][3] ) );
  DFEC1 \ram_reg[11][3]  ( .D(n199), .E(n226), .C(CLK), .RN(n164), .Q(
        \ram[11][3] ) );
  DFEC1 \ram_reg[13][3]  ( .D(n199), .E(n222), .C(CLK), .RN(n163), .Q(
        \ram[13][3] ) );
  DFEC1 \ram_reg[20][3]  ( .D(n198), .E(n243), .C(CLK), .RN(n160), .Q(
        \ram[20][3] ) );
  DFEC1 \ram_reg[25][3]  ( .D(n197), .E(n232), .C(CLK), .RN(n157), .Q(
        \ram[25][3] ) );
  DFEC1 \ram_reg[29][3]  ( .D(n197), .E(n224), .C(CLK), .RN(n155), .Q(
        \ram[29][3] ) );
  DFEC1 \ram_reg[31][3]  ( .D(n197), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][3] ) );
  DFEP1 \ram_reg[3][3]  ( .D(n200), .E(n225), .C(CLK), .SN(n174), .Q(
        \ram[3][3] ) );
  DFEP1 \ram_reg[4][3]  ( .D(n200), .E(n241), .C(CLK), .SN(n175), .Q(
        \ram[4][3] ) );
  DFEP1 \ram_reg[7][3]  ( .D(n200), .E(n217), .C(CLK), .SN(n178), .Q(
        \ram[7][3] ) );
  DFEP1 \ram_reg[8][3]  ( .D(n199), .E(n234), .C(CLK), .SN(n180), .Q(
        \ram[8][3] ) );
  DFEP1 \ram_reg[12][3]  ( .D(n199), .E(n242), .C(CLK), .SN(n171), .Q(
        \ram[12][3] ) );
  DFEP1 \ram_reg[15][3]  ( .D(n199), .E(n218), .C(CLK), .SN(n177), .Q(
        \ram[15][3] ) );
  DFEP1 \ram_reg[16][3]  ( .D(n198), .E(n235), .C(CLK), .SN(n181), .Q(
        \ram[16][3] ) );
  DFEP1 \ram_reg[17][3]  ( .D(n198), .E(n231), .C(CLK), .SN(n180), .Q(
        \ram[17][3] ) );
  DFEP1 \ram_reg[19][3]  ( .D(n198), .E(n227), .C(CLK), .SN(n179), .Q(
        \ram[19][3] ) );
  DFEP1 \ram_reg[21][3]  ( .D(n198), .E(n223), .C(CLK), .SN(n177), .Q(
        \ram[21][3] ) );
  DFEP1 \ram_reg[23][3]  ( .D(n198), .E(n219), .C(CLK), .SN(n176), .Q(
        \ram[23][3] ) );
  DFEP1 \ram_reg[24][3]  ( .D(n197), .E(n236), .C(CLK), .SN(n175), .Q(
        \ram[24][3] ) );
  DFEP1 \ram_reg[27][3]  ( .D(n197), .E(n228), .C(CLK), .SN(n173), .Q(
        \ram[27][3] ) );
  DFEP1 \ram_reg[28][3]  ( .D(n197), .E(n244), .C(CLK), .SN(n172), .Q(
        \ram[28][3] ) );
  DFEC1 \ram_reg[2][2]  ( .D(n196), .E(n237), .C(CLK), .RN(n166), .Q(
        \ram[2][2] ) );
  DFEC1 \ram_reg[2][1]  ( .D(n192), .E(n237), .C(CLK), .RN(n166), .Q(
        \ram[2][1] ) );
  DFEC1 \ram_reg[6][1]  ( .D(n192), .E(n245), .C(CLK), .RN(n168), .Q(
        \ram[6][1] ) );
  DFEC1 \ram_reg[10][1]  ( .D(n191), .E(n238), .C(CLK), .RN(n169), .Q(
        \ram[10][1] ) );
  DFEC1 \ram_reg[14][0]  ( .D(n187), .E(n246), .C(CLK), .RN(n162), .Q(
        \ram[14][0] ) );
  DFEC1 \ram_reg[18][1]  ( .D(n190), .E(n239), .C(CLK), .RN(n161), .Q(
        \ram[18][1] ) );
  DFEC1 \ram_reg[18][0]  ( .D(n186), .E(n239), .C(CLK), .RN(n161), .Q(
        \ram[18][0] ) );
  DFEC1 \ram_reg[22][2]  ( .D(n194), .E(n247), .C(CLK), .RN(n158), .Q(
        \ram[22][2] ) );
  DFEC1 \ram_reg[26][1]  ( .D(n189), .E(n240), .C(CLK), .RN(n156), .Q(
        \ram[26][1] ) );
  DFEC1 \ram_reg[26][0]  ( .D(n185), .E(n240), .C(CLK), .RN(n156), .Q(
        \ram[26][0] ) );
  DFEC1 \ram_reg[30][1]  ( .D(n189), .E(n248), .C(CLK), .RN(n155), .Q(
        \ram[30][1] ) );
  DFEC1 \ram_reg[30][0]  ( .D(n185), .E(n248), .C(CLK), .RN(n154), .Q(
        \ram[30][0] ) );
  DFEP1 \ram_reg[2][0]  ( .D(n188), .E(n237), .C(CLK), .SN(n172), .Q(
        \ram[2][0] ) );
  DFEP1 \ram_reg[6][2]  ( .D(n196), .E(n245), .C(CLK), .SN(n178), .Q(
        \ram[6][2] ) );
  DFEP1 \ram_reg[6][0]  ( .D(n188), .E(n245), .C(CLK), .SN(n178), .Q(
        \ram[6][0] ) );
  DFEP1 \ram_reg[10][2]  ( .D(n195), .E(n238), .C(CLK), .SN(n171), .Q(
        \ram[10][2] ) );
  DFEP1 \ram_reg[10][0]  ( .D(n187), .E(n238), .C(CLK), .SN(n170), .Q(
        \ram[10][0] ) );
  DFEP1 \ram_reg[14][2]  ( .D(n195), .E(n246), .C(CLK), .SN(n176), .Q(
        \ram[14][2] ) );
  DFEP1 \ram_reg[14][1]  ( .D(n191), .E(n246), .C(CLK), .SN(n177), .Q(
        \ram[14][1] ) );
  DFEP1 \ram_reg[18][2]  ( .D(n194), .E(n239), .C(CLK), .SN(n179), .Q(
        \ram[18][2] ) );
  DFEP1 \ram_reg[22][1]  ( .D(n190), .E(n247), .C(CLK), .SN(n176), .Q(
        \ram[22][1] ) );
  DFEP1 \ram_reg[22][0]  ( .D(n186), .E(n247), .C(CLK), .SN(n176), .Q(
        \ram[22][0] ) );
  DFEP1 \ram_reg[26][2]  ( .D(n193), .E(n240), .C(CLK), .SN(n174), .Q(
        \ram[26][2] ) );
  DFEP1 \ram_reg[30][2]  ( .D(n193), .E(n248), .C(CLK), .SN(n171), .Q(
        \ram[30][2] ) );
  DFEC1 \ram_reg[0][2]  ( .D(n196), .E(n233), .C(CLK), .RN(n164), .Q(
        \ram[0][2] ) );
  DFEC1 \ram_reg[0][1]  ( .D(n192), .E(n233), .C(CLK), .RN(n164), .Q(
        \ram[0][1] ) );
  DFEC1 \ram_reg[0][0]  ( .D(n188), .E(n233), .C(CLK), .RN(n164), .Q(
        \ram[0][0] ) );
  DFEC1 \ram_reg[1][1]  ( .D(n192), .E(n229), .C(CLK), .RN(n165), .Q(
        \ram[1][1] ) );
  DFEC1 \ram_reg[1][0]  ( .D(n188), .E(n229), .C(CLK), .RN(n165), .Q(
        \ram[1][0] ) );
  DFEC1 \ram_reg[3][1]  ( .D(n192), .E(n225), .C(CLK), .RN(n166), .Q(
        \ram[3][1] ) );
  DFEC1 \ram_reg[4][0]  ( .D(n188), .E(n241), .C(CLK), .RN(n166), .Q(
        \ram[4][0] ) );
  DFEC1 \ram_reg[5][1]  ( .D(n192), .E(n221), .C(CLK), .RN(n167), .Q(
        \ram[5][1] ) );
  DFEC1 \ram_reg[5][0]  ( .D(n188), .E(n221), .C(CLK), .RN(n167), .Q(
        \ram[5][0] ) );
  DFEC1 \ram_reg[7][1]  ( .D(n192), .E(n217), .C(CLK), .RN(n168), .Q(
        \ram[7][1] ) );
  DFEC1 \ram_reg[7][0]  ( .D(n188), .E(n217), .C(CLK), .RN(n168), .Q(
        \ram[7][0] ) );
  DFEC1 \ram_reg[8][2]  ( .D(n195), .E(n234), .C(CLK), .RN(n168), .Q(
        \ram[8][2] ) );
  DFEC1 \ram_reg[8][1]  ( .D(n191), .E(n234), .C(CLK), .RN(n168), .Q(
        \ram[8][1] ) );
  DFEC1 \ram_reg[8][0]  ( .D(n187), .E(n234), .C(CLK), .RN(n168), .Q(
        \ram[8][0] ) );
  DFEC1 \ram_reg[9][2]  ( .D(n195), .E(n230), .C(CLK), .RN(n170), .Q(
        \ram[9][2] ) );
  DFEC1 \ram_reg[11][2]  ( .D(n195), .E(n226), .C(CLK), .RN(n163), .Q(
        \ram[11][2] ) );
  DFEC1 \ram_reg[11][1]  ( .D(n191), .E(n226), .C(CLK), .RN(n163), .Q(
        \ram[11][1] ) );
  DFEC1 \ram_reg[12][2]  ( .D(n195), .E(n242), .C(CLK), .RN(n163), .Q(
        \ram[12][2] ) );
  DFEC1 \ram_reg[12][0]  ( .D(n187), .E(n242), .C(CLK), .RN(n163), .Q(
        \ram[12][0] ) );
  DFEC1 \ram_reg[13][1]  ( .D(n191), .E(n222), .C(CLK), .RN(n163), .Q(
        \ram[13][1] ) );
  DFEC1 \ram_reg[13][0]  ( .D(n187), .E(n222), .C(CLK), .RN(n163), .Q(
        \ram[13][0] ) );
  DFEC1 \ram_reg[15][2]  ( .D(n195), .E(n218), .C(CLK), .RN(n162), .Q(
        \ram[15][2] ) );
  DFEC1 \ram_reg[15][0]  ( .D(n187), .E(n218), .C(CLK), .RN(n164), .Q(
        \ram[15][0] ) );
  DFEC1 \ram_reg[16][2]  ( .D(n194), .E(n235), .C(CLK), .RN(n161), .Q(
        \ram[16][2] ) );
  DFEC1 \ram_reg[16][0]  ( .D(n186), .E(n235), .C(CLK), .RN(n161), .Q(
        \ram[16][0] ) );
  DFEC1 \ram_reg[17][0]  ( .D(n186), .E(n231), .C(CLK), .RN(n161), .Q(
        \ram[17][0] ) );
  DFEC1 \ram_reg[19][2]  ( .D(n194), .E(n227), .C(CLK), .RN(n160), .Q(
        \ram[19][2] ) );
  DFEC1 \ram_reg[19][0]  ( .D(n186), .E(n227), .C(CLK), .RN(n160), .Q(
        \ram[19][0] ) );
  DFEC1 \ram_reg[20][2]  ( .D(n194), .E(n243), .C(CLK), .RN(n160), .Q(
        \ram[20][2] ) );
  DFEC1 \ram_reg[20][1]  ( .D(n190), .E(n243), .C(CLK), .RN(n159), .Q(
        \ram[20][1] ) );
  DFEC1 \ram_reg[21][1]  ( .D(n190), .E(n223), .C(CLK), .RN(n159), .Q(
        \ram[21][1] ) );
  DFEC1 \ram_reg[23][2]  ( .D(n194), .E(n219), .C(CLK), .RN(n158), .Q(
        \ram[23][2] ) );
  DFEC1 \ram_reg[23][1]  ( .D(n190), .E(n219), .C(CLK), .RN(n158), .Q(
        \ram[23][1] ) );
  DFEC1 \ram_reg[23][0]  ( .D(n186), .E(n219), .C(CLK), .RN(n158), .Q(
        \ram[23][0] ) );
  DFEC1 \ram_reg[24][1]  ( .D(n189), .E(n236), .C(CLK), .RN(n158), .Q(
        \ram[24][1] ) );
  DFEC1 \ram_reg[24][0]  ( .D(n185), .E(n236), .C(CLK), .RN(n158), .Q(
        \ram[24][0] ) );
  DFEC1 \ram_reg[25][1]  ( .D(n189), .E(n232), .C(CLK), .RN(n157), .Q(
        \ram[25][1] ) );
  DFEC1 \ram_reg[27][0]  ( .D(n185), .E(n228), .C(CLK), .RN(n156), .Q(
        \ram[27][0] ) );
  DFEC1 \ram_reg[28][1]  ( .D(n189), .E(n244), .C(CLK), .RN(n156), .Q(
        \ram[28][1] ) );
  DFEC1 \ram_reg[29][2]  ( .D(n193), .E(n224), .C(CLK), .RN(n155), .Q(
        \ram[29][2] ) );
  DFEC1 \ram_reg[29][1]  ( .D(n189), .E(n224), .C(CLK), .RN(n155), .Q(
        \ram[29][1] ) );
  DFEC1 \ram_reg[31][2]  ( .D(n193), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][2] ) );
  DFEC1 \ram_reg[31][1]  ( .D(n189), .E(n220), .C(CLK), .RN(n154), .Q(
        \ram[31][1] ) );
  DFEC1 \ram_reg[31][0]  ( .D(n185), .E(n220), .C(CLK), .RN(n162), .Q(
        \ram[31][0] ) );
  DFEP1 \ram_reg[1][2]  ( .D(n196), .E(n229), .C(CLK), .SN(n170), .Q(
        \ram[1][2] ) );
  DFEP1 \ram_reg[3][2]  ( .D(n196), .E(n225), .C(CLK), .SN(n174), .Q(
        \ram[3][2] ) );
  DFEP1 \ram_reg[3][0]  ( .D(n188), .E(n225), .C(CLK), .SN(n174), .Q(
        \ram[3][0] ) );
  DFEP1 \ram_reg[4][2]  ( .D(n196), .E(n241), .C(CLK), .SN(n175), .Q(
        \ram[4][2] ) );
  DFEP1 \ram_reg[4][1]  ( .D(n192), .E(n241), .C(CLK), .SN(n175), .Q(
        \ram[4][1] ) );
  DFEP1 \ram_reg[5][2]  ( .D(n196), .E(n221), .C(CLK), .SN(n177), .Q(
        \ram[5][2] ) );
  DFEP1 \ram_reg[7][2]  ( .D(n196), .E(n217), .C(CLK), .SN(n178), .Q(
        \ram[7][2] ) );
  DFEP1 \ram_reg[9][1]  ( .D(n191), .E(n230), .C(CLK), .SN(n177), .Q(
        \ram[9][1] ) );
  DFEP1 \ram_reg[9][0]  ( .D(n187), .E(n230), .C(CLK), .SN(n177), .Q(
        \ram[9][0] ) );
  DFEP1 \ram_reg[11][0]  ( .D(n187), .E(n226), .C(CLK), .SN(n170), .Q(
        \ram[11][0] ) );
  DFEP1 \ram_reg[12][1]  ( .D(n191), .E(n242), .C(CLK), .SN(n170), .Q(
        \ram[12][1] ) );
  DFEP1 \ram_reg[13][2]  ( .D(n195), .E(n222), .C(CLK), .SN(n172), .Q(
        \ram[13][2] ) );
  DFEP1 \ram_reg[15][1]  ( .D(n191), .E(n218), .C(CLK), .SN(n178), .Q(
        \ram[15][1] ) );
  DFEP1 \ram_reg[16][1]  ( .D(n190), .E(n235), .C(CLK), .SN(n170), .Q(
        \ram[16][1] ) );
  DFEP1 \ram_reg[17][2]  ( .D(n194), .E(n231), .C(CLK), .SN(n180), .Q(
        \ram[17][2] ) );
  DFEP1 \ram_reg[17][1]  ( .D(n190), .E(n231), .C(CLK), .SN(n180), .Q(
        \ram[17][1] ) );
  DFEP1 \ram_reg[19][1]  ( .D(n190), .E(n227), .C(CLK), .SN(n179), .Q(
        \ram[19][1] ) );
  DFEP1 \ram_reg[20][0]  ( .D(n186), .E(n243), .C(CLK), .SN(n178), .Q(
        \ram[20][0] ) );
  DFEP1 \ram_reg[21][2]  ( .D(n194), .E(n223), .C(CLK), .SN(n177), .Q(
        \ram[21][2] ) );
  DFEP1 \ram_reg[21][0]  ( .D(n186), .E(n223), .C(CLK), .SN(n177), .Q(
        \ram[21][0] ) );
  DFEP1 \ram_reg[24][2]  ( .D(n193), .E(n236), .C(CLK), .SN(n175), .Q(
        \ram[24][2] ) );
  DFEP1 \ram_reg[25][2]  ( .D(n193), .E(n232), .C(CLK), .SN(n174), .Q(
        \ram[25][2] ) );
  DFEP1 \ram_reg[25][0]  ( .D(n185), .E(n232), .C(CLK), .SN(n174), .Q(
        \ram[25][0] ) );
  DFEP1 \ram_reg[27][2]  ( .D(n193), .E(n228), .C(CLK), .SN(n172), .Q(
        \ram[27][2] ) );
  DFEP1 \ram_reg[27][1]  ( .D(n189), .E(n228), .C(CLK), .SN(n173), .Q(
        \ram[27][1] ) );
  DFEP1 \ram_reg[28][2]  ( .D(n193), .E(n244), .C(CLK), .SN(n172), .Q(
        \ram[28][2] ) );
  DFEP1 \ram_reg[28][0]  ( .D(n185), .E(n244), .C(CLK), .SN(n171), .Q(
        \ram[28][0] ) );
  DFEP1 \ram_reg[29][0]  ( .D(n185), .E(n224), .C(CLK), .SN(n171), .Q(
        \ram[29][0] ) );
  NOR31 U2 ( .A(n139), .B(wb), .C(n250), .Q(n40) );
  BUF2 U3 ( .A(N11), .Q(n125) );
  BUF2 U4 ( .A(n132), .Q(n127) );
  BUF2 U5 ( .A(n132), .Q(n126) );
  BUF2 U6 ( .A(n133), .Q(n128) );
  BUF2 U7 ( .A(n133), .Q(n129) );
  BUF2 U8 ( .A(n134), .Q(n130) );
  BUF2 U9 ( .A(n134), .Q(n131) );
  BUF2 U10 ( .A(n182), .Q(n136) );
  BUF2 U11 ( .A(n182), .Q(n137) );
  BUF2 U12 ( .A(n182), .Q(n135) );
  BUF2 U13 ( .A(N11), .Q(n132) );
  BUF2 U14 ( .A(n182), .Q(n138) );
  BUF2 U15 ( .A(N11), .Q(n133) );
  BUF2 U16 ( .A(N11), .Q(n134) );
  INV3 U17 ( .A(n183), .Q(n182) );
  NOR31 U18 ( .A(n184), .B(n183), .C(n249), .Q(n41) );
  NOR31 U19 ( .A(n184), .B(n182), .C(n249), .Q(n43) );
  NOR31 U20 ( .A(n183), .B(N11), .C(n249), .Q(n45) );
  NOR31 U21 ( .A(n182), .B(N11), .C(n249), .Q(n47) );
  BUF2 U22 ( .A(n148), .Q(n170) );
  BUF2 U23 ( .A(n151), .Q(n176) );
  BUF2 U24 ( .A(n148), .Q(n171) );
  BUF2 U25 ( .A(n153), .Q(n180) );
  BUF2 U26 ( .A(n152), .Q(n179) );
  BUF2 U27 ( .A(n152), .Q(n178) );
  BUF2 U28 ( .A(n151), .Q(n177) );
  BUF2 U29 ( .A(n150), .Q(n175) );
  BUF2 U30 ( .A(n150), .Q(n174) );
  BUF2 U31 ( .A(n149), .Q(n173) );
  BUF2 U32 ( .A(n149), .Q(n172) );
  BUF2 U33 ( .A(n140), .Q(n155) );
  BUF2 U34 ( .A(n141), .Q(n156) );
  BUF2 U35 ( .A(n141), .Q(n157) );
  BUF2 U36 ( .A(n142), .Q(n158) );
  BUF2 U37 ( .A(n142), .Q(n159) );
  BUF2 U38 ( .A(n143), .Q(n160) );
  BUF2 U39 ( .A(n143), .Q(n161) );
  BUF2 U40 ( .A(n144), .Q(n162) );
  BUF2 U41 ( .A(n144), .Q(n163) );
  BUF2 U42 ( .A(n147), .Q(n169) );
  BUF2 U43 ( .A(n146), .Q(n167) );
  BUF2 U44 ( .A(n147), .Q(n168) );
  BUF2 U45 ( .A(n145), .Q(n165) );
  BUF2 U46 ( .A(n145), .Q(n164) );
  BUF2 U47 ( .A(n146), .Q(n166) );
  BUF2 U48 ( .A(n140), .Q(n154) );
  BUF2 U49 ( .A(n153), .Q(n181) );
  INV3 U50 ( .A(N10), .Q(n183) );
  INV3 U51 ( .A(N11), .Q(n184) );
  INV3 U52 ( .A(N13), .Q(n139) );
  INV3 U53 ( .A(n39), .Q(n220) );
  NAND22 U54 ( .A(n40), .B(n41), .Q(n39) );
  INV3 U55 ( .A(n82), .Q(n233) );
  NAND22 U56 ( .A(n75), .B(n55), .Q(n82) );
  INV3 U57 ( .A(n42), .Q(n248) );
  NAND22 U58 ( .A(n43), .B(n40), .Q(n42) );
  INV3 U59 ( .A(n44), .Q(n224) );
  NAND22 U60 ( .A(n45), .B(n40), .Q(n44) );
  INV3 U61 ( .A(n50), .Q(n240) );
  NAND22 U62 ( .A(n51), .B(n40), .Q(n50) );
  INV3 U63 ( .A(n70), .Q(n226) );
  NAND22 U64 ( .A(n66), .B(n49), .Q(n70) );
  INV3 U65 ( .A(n77), .Q(n221) );
  NAND22 U66 ( .A(n75), .B(n45), .Q(n77) );
  INV3 U67 ( .A(n80), .Q(n237) );
  NAND22 U68 ( .A(n75), .B(n51), .Q(n80) );
  INV3 U69 ( .A(n81), .Q(n229) );
  NAND22 U70 ( .A(n75), .B(n53), .Q(n81) );
  INV3 U71 ( .A(n60), .Q(n243) );
  NAND22 U72 ( .A(n57), .B(n47), .Q(n60) );
  INV3 U73 ( .A(n52), .Q(n232) );
  NAND22 U74 ( .A(n53), .B(n40), .Q(n52) );
  INV3 U75 ( .A(n72), .Q(n230) );
  NAND22 U76 ( .A(n66), .B(n53), .Q(n72) );
  INV3 U77 ( .A(n76), .Q(n245) );
  NAND22 U78 ( .A(n75), .B(n43), .Q(n76) );
  INV3 U79 ( .A(n58), .Q(n247) );
  NAND22 U80 ( .A(n57), .B(n43), .Q(n58) );
  INV3 U81 ( .A(n71), .Q(n238) );
  NAND22 U82 ( .A(n66), .B(n51), .Q(n71) );
  INV3 U83 ( .A(n59), .Q(n223) );
  NAND22 U84 ( .A(n57), .B(n45), .Q(n59) );
  INV3 U85 ( .A(n65), .Q(n218) );
  NAND22 U86 ( .A(n66), .B(n41), .Q(n65) );
  INV3 U87 ( .A(n67), .Q(n246) );
  NAND22 U88 ( .A(n66), .B(n43), .Q(n67) );
  INV3 U89 ( .A(n63), .Q(n231) );
  NAND22 U90 ( .A(n57), .B(n53), .Q(n63) );
  INV3 U91 ( .A(n64), .Q(n235) );
  NAND22 U92 ( .A(n57), .B(n55), .Q(n64) );
  INV3 U93 ( .A(n68), .Q(n222) );
  NAND22 U94 ( .A(n66), .B(n45), .Q(n68) );
  INV3 U95 ( .A(n69), .Q(n242) );
  NAND22 U96 ( .A(n66), .B(n47), .Q(n69) );
  INV3 U97 ( .A(n73), .Q(n234) );
  NAND22 U98 ( .A(n66), .B(n55), .Q(n73) );
  INV3 U99 ( .A(n56), .Q(n219) );
  NAND22 U100 ( .A(n57), .B(n41), .Q(n56) );
  INV3 U101 ( .A(n61), .Q(n227) );
  NAND22 U102 ( .A(n57), .B(n49), .Q(n61) );
  INV3 U103 ( .A(n62), .Q(n239) );
  NAND22 U104 ( .A(n57), .B(n51), .Q(n62) );
  INV3 U105 ( .A(n54), .Q(n236) );
  NAND22 U106 ( .A(n55), .B(n40), .Q(n54) );
  INV3 U107 ( .A(n74), .Q(n217) );
  NAND22 U108 ( .A(n75), .B(n41), .Q(n74) );
  INV3 U109 ( .A(n46), .Q(n244) );
  NAND22 U110 ( .A(n47), .B(n40), .Q(n46) );
  INV3 U111 ( .A(n48), .Q(n228) );
  NAND22 U112 ( .A(n49), .B(n40), .Q(n48) );
  INV3 U113 ( .A(n78), .Q(n241) );
  NAND22 U114 ( .A(n75), .B(n47), .Q(n78) );
  INV3 U115 ( .A(n79), .Q(n225) );
  NAND22 U116 ( .A(n75), .B(n49), .Q(n79) );
  INV3 U117 ( .A(N14), .Q(n250) );
  NOR31 U118 ( .A(n183), .B(N12), .C(n184), .Q(n49) );
  NOR31 U119 ( .A(n182), .B(N12), .C(n184), .Q(n51) );
  NOR31 U120 ( .A(N11), .B(N12), .C(n183), .Q(n53) );
  NOR31 U121 ( .A(N11), .B(N12), .C(n182), .Q(n55) );
  INV3 U122 ( .A(N12), .Q(n249) );
  BUF2 U123 ( .A(n251), .Q(n141) );
  BUF2 U124 ( .A(n251), .Q(n142) );
  BUF2 U125 ( .A(n251), .Q(n143) );
  BUF2 U126 ( .A(n251), .Q(n144) );
  BUF2 U127 ( .A(n251), .Q(n153) );
  BUF2 U128 ( .A(n251), .Q(n152) );
  BUF2 U129 ( .A(n251), .Q(n151) );
  BUF2 U130 ( .A(n251), .Q(n150) );
  BUF2 U131 ( .A(n251), .Q(n149) );
  BUF2 U132 ( .A(n251), .Q(n147) );
  BUF2 U133 ( .A(n251), .Q(n148) );
  BUF2 U134 ( .A(n251), .Q(n145) );
  BUF2 U135 ( .A(n251), .Q(n146) );
  BUF2 U136 ( .A(n251), .Q(n140) );
  IMUX40 U137 ( .A(\ram[28][1] ), .B(\ram[29][1] ), .C(\ram[30][1] ), .D(
        \ram[31][1] ), .S0(n136), .S1(n125), .Q(n15) );
  IMUX40 U138 ( .A(\ram[16][1] ), .B(\ram[17][1] ), .C(\ram[18][1] ), .D(
        \ram[19][1] ), .S0(n136), .S1(n126), .Q(n12) );
  IMUX40 U139 ( .A(\ram[24][1] ), .B(\ram[25][1] ), .C(\ram[26][1] ), .D(
        \ram[27][1] ), .S0(n136), .S1(n125), .Q(n13) );
  IMUX40 U140 ( .A(\ram[12][1] ), .B(\ram[13][1] ), .C(\ram[14][1] ), .D(
        \ram[15][1] ), .S0(n136), .S1(n126), .Q(n20) );
  IMUX40 U141 ( .A(\ram[0][1] ), .B(\ram[1][1] ), .C(\ram[2][1] ), .D(
        \ram[3][1] ), .S0(n136), .S1(n126), .Q(n17) );
  IMUX40 U142 ( .A(\ram[8][1] ), .B(\ram[9][1] ), .C(\ram[10][1] ), .D(
        \ram[11][1] ), .S0(n136), .S1(n126), .Q(n18) );
  IMUX40 U143 ( .A(\ram[20][1] ), .B(\ram[21][1] ), .C(\ram[22][1] ), .D(
        \ram[23][1] ), .S0(n136), .S1(n126), .Q(n14) );
  MUX22 U144 ( .A(n16), .B(n11), .S(N14), .Q(data_out[1]) );
  IMUX40 U145 ( .A(n17), .B(n18), .C(n19), .D(n20), .S0(N13), .S1(N12), .Q(n16) );
  IMUX40 U146 ( .A(n12), .B(n13), .C(n14), .D(n15), .S0(N13), .S1(N12), .Q(n11) );
  IMUX40 U147 ( .A(\ram[4][1] ), .B(\ram[5][1] ), .C(\ram[6][1] ), .D(
        \ram[7][1] ), .S0(n136), .S1(n126), .Q(n19) );
  IMUX40 U148 ( .A(\ram[12][0] ), .B(\ram[13][0] ), .C(\ram[14][0] ), .D(
        \ram[15][0] ), .S0(n136), .S1(n125), .Q(n10) );
  IMUX40 U149 ( .A(\ram[0][0] ), .B(\ram[1][0] ), .C(\ram[2][0] ), .D(
        \ram[3][0] ), .S0(n136), .S1(n125), .Q(n7) );
  IMUX40 U150 ( .A(\ram[8][0] ), .B(\ram[9][0] ), .C(\ram[10][0] ), .D(
        \ram[11][0] ), .S0(n136), .S1(n125), .Q(n8) );
  IMUX40 U151 ( .A(\ram[28][2] ), .B(\ram[29][2] ), .C(\ram[30][2] ), .D(
        \ram[31][2] ), .S0(n137), .S1(n126), .Q(n25) );
  IMUX40 U152 ( .A(\ram[16][2] ), .B(\ram[17][2] ), .C(\ram[18][2] ), .D(
        \ram[19][2] ), .S0(n137), .S1(n127), .Q(n22) );
  IMUX40 U153 ( .A(\ram[24][2] ), .B(\ram[25][2] ), .C(\ram[26][2] ), .D(
        \ram[27][2] ), .S0(n137), .S1(n126), .Q(n23) );
  IMUX40 U154 ( .A(\ram[12][2] ), .B(\ram[13][2] ), .C(\ram[14][2] ), .D(
        \ram[15][2] ), .S0(n137), .S1(n127), .Q(n30) );
  IMUX40 U155 ( .A(\ram[0][2] ), .B(\ram[1][2] ), .C(\ram[2][2] ), .D(
        \ram[3][2] ), .S0(n137), .S1(n127), .Q(n27) );
  IMUX40 U156 ( .A(\ram[8][2] ), .B(\ram[9][2] ), .C(\ram[10][2] ), .D(
        \ram[11][2] ), .S0(n137), .S1(n127), .Q(n28) );
  IMUX40 U157 ( .A(\ram[28][3] ), .B(\ram[29][3] ), .C(\ram[30][3] ), .D(
        \ram[31][3] ), .S0(n137), .S1(n127), .Q(n35) );
  IMUX40 U158 ( .A(\ram[16][3] ), .B(\ram[17][3] ), .C(\ram[18][3] ), .D(
        \ram[19][3] ), .S0(n137), .S1(n127), .Q(n32) );
  IMUX40 U159 ( .A(\ram[24][3] ), .B(\ram[25][3] ), .C(\ram[26][3] ), .D(
        \ram[27][3] ), .S0(n137), .S1(n127), .Q(n33) );
  IMUX40 U160 ( .A(\ram[30][0] ), .B(\ram[31][0] ), .C(\ram[28][0] ), .D(
        \ram[29][0] ), .S0(n135), .S1(n184), .Q(n5) );
  IMUX40 U161 ( .A(\ram[16][0] ), .B(\ram[17][0] ), .C(\ram[18][0] ), .D(
        \ram[19][0] ), .S0(n135), .S1(n125), .Q(n2) );
  IMUX40 U162 ( .A(\ram[24][0] ), .B(\ram[25][0] ), .C(\ram[26][0] ), .D(
        \ram[27][0] ), .S0(n135), .S1(n125), .Q(n3) );
  IMUX40 U163 ( .A(\ram[4][0] ), .B(\ram[5][0] ), .C(\ram[6][0] ), .D(
        \ram[7][0] ), .S0(n136), .S1(n125), .Q(n9) );
  IMUX40 U164 ( .A(\ram[20][2] ), .B(\ram[21][2] ), .C(\ram[22][2] ), .D(
        \ram[23][2] ), .S0(n137), .S1(n126), .Q(n24) );
  MUX22 U165 ( .A(n6), .B(n1), .S(N14), .Q(data_out[0]) );
  IMUX40 U166 ( .A(n2), .B(n3), .C(n4), .D(n5), .S0(N13), .S1(N12), .Q(n1) );
  IMUX40 U167 ( .A(n7), .B(n8), .C(n9), .D(n10), .S0(N13), .S1(N12), .Q(n6) );
  IMUX40 U168 ( .A(\ram[20][0] ), .B(\ram[21][0] ), .C(\ram[22][0] ), .D(
        \ram[23][0] ), .S0(n135), .S1(n125), .Q(n4) );
  MUX22 U169 ( .A(n26), .B(n21), .S(N14), .Q(data_out[2]) );
  IMUX40 U170 ( .A(n27), .B(n28), .C(n29), .D(n30), .S0(N13), .S1(N12), .Q(n26) );
  IMUX40 U171 ( .A(n22), .B(n23), .C(n24), .D(n25), .S0(N13), .S1(N12), .Q(n21) );
  IMUX40 U172 ( .A(\ram[4][2] ), .B(\ram[5][2] ), .C(\ram[6][2] ), .D(
        \ram[7][2] ), .S0(n137), .S1(n127), .Q(n29) );
  MUX22 U173 ( .A(n36), .B(n31), .S(N14), .Q(data_out[3]) );
  IMUX40 U174 ( .A(n37), .B(n38), .C(n83), .D(n84), .S0(N13), .S1(N12), .Q(n36) );
  IMUX40 U175 ( .A(n32), .B(n33), .C(n34), .D(n35), .S0(N13), .S1(N12), .Q(n31) );
  IMUX40 U176 ( .A(\ram[4][3] ), .B(\ram[5][3] ), .C(\ram[6][3] ), .D(
        \ram[7][3] ), .S0(n138), .S1(n128), .Q(n83) );
  IMUX40 U177 ( .A(\ram[12][3] ), .B(\ram[13][3] ), .C(\ram[14][3] ), .D(
        \ram[15][3] ), .S0(n138), .S1(n128), .Q(n84) );
  IMUX40 U178 ( .A(\ram[0][3] ), .B(\ram[1][3] ), .C(\ram[2][3] ), .D(
        \ram[3][3] ), .S0(n138), .S1(n128), .Q(n37) );
  IMUX40 U179 ( .A(\ram[8][3] ), .B(\ram[9][3] ), .C(\ram[10][3] ), .D(
        \ram[11][3] ), .S0(n138), .S1(n128), .Q(n38) );
  IMUX40 U180 ( .A(\ram[28][4] ), .B(\ram[29][4] ), .C(\ram[30][4] ), .D(
        \ram[31][4] ), .S0(n138), .S1(n128), .Q(n89) );
  IMUX40 U181 ( .A(\ram[16][4] ), .B(\ram[17][4] ), .C(\ram[18][4] ), .D(
        \ram[19][4] ), .S0(n138), .S1(n128), .Q(n86) );
  IMUX40 U182 ( .A(\ram[24][4] ), .B(\ram[25][4] ), .C(\ram[26][4] ), .D(
        \ram[27][4] ), .S0(n138), .S1(n128), .Q(n87) );
  IMUX40 U183 ( .A(\ram[12][4] ), .B(\ram[13][4] ), .C(\ram[14][4] ), .D(
        \ram[15][4] ), .S0(n138), .S1(n128), .Q(n94) );
  IMUX40 U184 ( .A(\ram[0][4] ), .B(\ram[1][4] ), .C(\ram[2][4] ), .D(
        \ram[3][4] ), .S0(n138), .S1(n129), .Q(n91) );
  IMUX40 U185 ( .A(\ram[8][4] ), .B(\ram[9][4] ), .C(\ram[10][4] ), .D(
        \ram[11][4] ), .S0(n138), .S1(n129), .Q(n92) );
  IMUX40 U186 ( .A(\ram[20][3] ), .B(\ram[21][3] ), .C(\ram[22][3] ), .D(
        \ram[23][3] ), .S0(n137), .S1(n127), .Q(n34) );
  IMUX40 U187 ( .A(\ram[20][4] ), .B(\ram[21][4] ), .C(\ram[22][4] ), .D(
        \ram[23][4] ), .S0(n138), .S1(n128), .Q(n88) );
  MUX22 U188 ( .A(n90), .B(n85), .S(N14), .Q(data_out[4]) );
  IMUX40 U189 ( .A(n91), .B(n92), .C(n93), .D(n94), .S0(N13), .S1(N12), .Q(n90) );
  IMUX40 U190 ( .A(n86), .B(n87), .C(n88), .D(n89), .S0(N13), .S1(N12), .Q(n85) );
  IMUX40 U191 ( .A(\ram[4][4] ), .B(\ram[5][4] ), .C(\ram[6][4] ), .D(
        \ram[7][4] ), .S0(n138), .S1(n129), .Q(n93) );
  IMUX40 U192 ( .A(\ram[28][5] ), .B(\ram[29][5] ), .C(\ram[30][5] ), .D(
        \ram[31][5] ), .S0(n138), .S1(n129), .Q(n99) );
  IMUX40 U193 ( .A(\ram[16][5] ), .B(\ram[17][5] ), .C(\ram[18][5] ), .D(
        \ram[19][5] ), .S0(n138), .S1(n129), .Q(n96) );
  IMUX40 U194 ( .A(\ram[24][5] ), .B(\ram[25][5] ), .C(\ram[26][5] ), .D(
        \ram[27][5] ), .S0(n138), .S1(n129), .Q(n97) );
  IMUX40 U195 ( .A(\ram[12][5] ), .B(\ram[13][5] ), .C(\ram[14][5] ), .D(
        \ram[15][5] ), .S0(n135), .S1(n129), .Q(n104) );
  IMUX40 U196 ( .A(\ram[0][5] ), .B(\ram[1][5] ), .C(\ram[2][5] ), .D(
        \ram[3][5] ), .S0(n135), .S1(n130), .Q(n101) );
  IMUX40 U197 ( .A(\ram[8][5] ), .B(\ram[9][5] ), .C(\ram[10][5] ), .D(
        \ram[11][5] ), .S0(n138), .S1(n129), .Q(n102) );
  IMUX40 U198 ( .A(\ram[28][6] ), .B(\ram[29][6] ), .C(\ram[30][6] ), .D(
        \ram[31][6] ), .S0(n138), .S1(n130), .Q(n109) );
  IMUX40 U199 ( .A(\ram[16][6] ), .B(\ram[17][6] ), .C(\ram[18][6] ), .D(
        \ram[19][6] ), .S0(n137), .S1(n130), .Q(n106) );
  IMUX40 U200 ( .A(\ram[24][6] ), .B(\ram[25][6] ), .C(\ram[26][6] ), .D(
        \ram[27][6] ), .S0(n137), .S1(n130), .Q(n107) );
  IMUX40 U201 ( .A(\ram[12][6] ), .B(\ram[13][6] ), .C(\ram[14][6] ), .D(
        \ram[15][6] ), .S0(n135), .S1(n130), .Q(n114) );
  IMUX40 U202 ( .A(\ram[0][6] ), .B(\ram[1][6] ), .C(\ram[2][6] ), .D(
        \ram[3][6] ), .S0(n135), .S1(n131), .Q(n111) );
  IMUX40 U203 ( .A(\ram[8][6] ), .B(\ram[9][6] ), .C(\ram[10][6] ), .D(
        \ram[11][6] ), .S0(n135), .S1(n130), .Q(n112) );
  IMUX40 U204 ( .A(\ram[20][5] ), .B(\ram[21][5] ), .C(\ram[22][5] ), .D(
        \ram[23][5] ), .S0(n135), .S1(n129), .Q(n98) );
  IMUX40 U205 ( .A(\ram[20][6] ), .B(\ram[21][6] ), .C(\ram[22][6] ), .D(
        \ram[23][6] ), .S0(n138), .S1(n130), .Q(n108) );
  MUX22 U206 ( .A(n100), .B(n95), .S(N14), .Q(data_out[5]) );
  IMUX40 U207 ( .A(n101), .B(n102), .C(n103), .D(n104), .S0(N13), .S1(N12), 
        .Q(n100) );
  IMUX40 U208 ( .A(n96), .B(n97), .C(n98), .D(n99), .S0(N13), .S1(N12), .Q(n95) );
  IMUX40 U209 ( .A(\ram[4][5] ), .B(\ram[5][5] ), .C(\ram[6][5] ), .D(
        \ram[7][5] ), .S0(n135), .S1(n130), .Q(n103) );
  MUX22 U210 ( .A(n110), .B(n105), .S(N14), .Q(data_out[6]) );
  IMUX40 U211 ( .A(n111), .B(n112), .C(n113), .D(n114), .S0(N13), .S1(N12), 
        .Q(n110) );
  IMUX40 U212 ( .A(n106), .B(n107), .C(n108), .D(n109), .S0(N13), .S1(N12), 
        .Q(n105) );
  IMUX40 U213 ( .A(\ram[4][6] ), .B(\ram[5][6] ), .C(\ram[6][6] ), .D(
        \ram[7][6] ), .S0(n137), .S1(n130), .Q(n113) );
  IMUX40 U214 ( .A(\ram[28][7] ), .B(\ram[29][7] ), .C(\ram[30][7] ), .D(
        \ram[31][7] ), .S0(n137), .S1(n131), .Q(n119) );
  IMUX40 U215 ( .A(\ram[16][7] ), .B(\ram[17][7] ), .C(\ram[18][7] ), .D(
        \ram[19][7] ), .S0(n138), .S1(n131), .Q(n116) );
  IMUX40 U216 ( .A(\ram[24][7] ), .B(\ram[25][7] ), .C(\ram[26][7] ), .D(
        \ram[27][7] ), .S0(n138), .S1(n131), .Q(n117) );
  IMUX40 U217 ( .A(\ram[12][7] ), .B(\ram[13][7] ), .C(\ram[14][7] ), .D(
        \ram[15][7] ), .S0(n135), .S1(n131), .Q(n124) );
  IMUX40 U218 ( .A(\ram[0][7] ), .B(\ram[1][7] ), .C(\ram[2][7] ), .D(
        \ram[3][7] ), .S0(n135), .S1(n131), .Q(n121) );
  IMUX40 U219 ( .A(\ram[8][7] ), .B(\ram[9][7] ), .C(\ram[10][7] ), .D(
        \ram[11][7] ), .S0(n135), .S1(n131), .Q(n122) );
  IMUX40 U220 ( .A(\ram[20][7] ), .B(\ram[21][7] ), .C(\ram[22][7] ), .D(
        \ram[23][7] ), .S0(n135), .S1(n131), .Q(n118) );
  MUX22 U221 ( .A(n120), .B(n115), .S(N14), .Q(data_out[7]) );
  IMUX40 U222 ( .A(n121), .B(n122), .C(n123), .D(n124), .S0(N13), .S1(N12), 
        .Q(n120) );
  IMUX40 U223 ( .A(n116), .B(n117), .C(n118), .D(n119), .S0(N13), .S1(N12), 
        .Q(n115) );
  IMUX40 U224 ( .A(\ram[4][7] ), .B(\ram[5][7] ), .C(\ram[6][7] ), .D(
        \ram[7][7] ), .S0(n135), .S1(n131), .Q(n123) );
  NOR31 U225 ( .A(N14), .B(wb), .C(n139), .Q(n66) );
  NOR31 U226 ( .A(N14), .B(wb), .C(N13), .Q(n75) );
  NOR31 U227 ( .A(N13), .B(wb), .C(n250), .Q(n57) );
  INV3 U228 ( .A(RESET), .Q(n251) );
  BUF2 U229 ( .A(data_in[0]), .Q(n185) );
  BUF2 U230 ( .A(data_in[1]), .Q(n189) );
  BUF2 U231 ( .A(data_in[2]), .Q(n193) );
  BUF2 U232 ( .A(data_in[3]), .Q(n197) );
  BUF2 U233 ( .A(data_in[4]), .Q(n201) );
  BUF2 U234 ( .A(data_in[5]), .Q(n205) );
  BUF2 U235 ( .A(data_in[6]), .Q(n209) );
  BUF2 U236 ( .A(data_in[7]), .Q(n213) );
  BUF2 U237 ( .A(data_in[0]), .Q(n186) );
  BUF2 U238 ( .A(data_in[1]), .Q(n190) );
  BUF2 U239 ( .A(data_in[2]), .Q(n194) );
  BUF2 U240 ( .A(data_in[3]), .Q(n198) );
  BUF2 U241 ( .A(data_in[4]), .Q(n202) );
  BUF2 U242 ( .A(data_in[5]), .Q(n206) );
  BUF2 U243 ( .A(data_in[6]), .Q(n210) );
  BUF2 U244 ( .A(data_in[7]), .Q(n214) );
  BUF2 U245 ( .A(data_in[0]), .Q(n187) );
  BUF2 U246 ( .A(data_in[1]), .Q(n191) );
  BUF2 U247 ( .A(data_in[2]), .Q(n195) );
  BUF2 U248 ( .A(data_in[3]), .Q(n199) );
  BUF2 U249 ( .A(data_in[4]), .Q(n203) );
  BUF2 U250 ( .A(data_in[5]), .Q(n207) );
  BUF2 U251 ( .A(data_in[6]), .Q(n211) );
  BUF2 U252 ( .A(data_in[7]), .Q(n215) );
  BUF2 U253 ( .A(data_in[0]), .Q(n188) );
  BUF2 U254 ( .A(data_in[1]), .Q(n192) );
  BUF2 U255 ( .A(data_in[2]), .Q(n196) );
  BUF2 U256 ( .A(data_in[3]), .Q(n200) );
  BUF2 U257 ( .A(data_in[4]), .Q(n204) );
  BUF2 U258 ( .A(data_in[5]), .Q(n208) );
  BUF2 U259 ( .A(data_in[6]), .Q(n212) );
  BUF2 U260 ( .A(data_in[7]), .Q(n216) );
endmodule


module MULT_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34;
  assign \A[5]  = A[5];
  assign SUM[5] = \A[5] ;
  assign \A[4]  = A[4];
  assign SUM[4] = \A[4] ;
  assign \A[3]  = A[3];
  assign SUM[3] = \A[3] ;
  assign \A[2]  = A[2];
  assign SUM[2] = \A[2] ;
  assign \A[1]  = A[1];
  assign SUM[1] = \A[1] ;
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  INV3 U2 ( .A(n26), .Q(n4) );
  INV3 U3 ( .A(n13), .Q(n5) );
  INV3 U4 ( .A(n14), .Q(n8) );
  INV3 U5 ( .A(n30), .Q(n6) );
  INV3 U6 ( .A(n25), .Q(n7) );
  INV3 U7 ( .A(n22), .Q(n2) );
  INV3 U8 ( .A(n28), .Q(n3) );
  INV3 U9 ( .A(n21), .Q(n1) );
  INV3 U10 ( .A(A[6]), .Q(n9) );
  INV3 U11 ( .A(B[6]), .Q(n10) );
  XNR20 U12 ( .A(n11), .B(n12), .Q(SUM[9]) );
  NAND20 U13 ( .A(n7), .B(n13), .Q(n12) );
  OAI210 U14 ( .A(n14), .B(n15), .C(n16), .Q(SUM[8]) );
  IMUX20 U15 ( .A(n17), .B(n18), .S(B[8]), .Q(n16) );
  NOR20 U16 ( .A(A[8]), .B(n8), .Q(n18) );
  XNR20 U17 ( .A(A[8]), .B(n14), .Q(n17) );
  XOR30 U18 ( .A(A[7]), .B(B[7]), .C(n19), .Q(SUM[7]) );
  AOI210 U19 ( .A(n10), .B(n9), .C(n19), .Q(SUM[6]) );
  XNR30 U20 ( .A(B[13]), .B(A[13]), .C(n20), .Q(SUM[13]) );
  AOI210 U21 ( .A(n2), .B(A[12]), .C(n1), .Q(n20) );
  OAI210 U22 ( .A(A[12]), .B(n2), .C(B[12]), .Q(n21) );
  XOR30 U23 ( .A(B[12]), .B(A[12]), .C(n2), .Q(SUM[12]) );
  AOI2110 U24 ( .A(n23), .B(A[11]), .C(n3), .D(n24), .Q(n22) );
  NOR40 U25 ( .A(n25), .B(n14), .C(n26), .D(n27), .Q(n24) );
  OAI220 U26 ( .A(A[11]), .B(B[11]), .C(A[8]), .D(B[8]), .Q(n27) );
  OAI210 U27 ( .A(A[11]), .B(n23), .C(B[11]), .Q(n28) );
  OAI210 U28 ( .A(n26), .B(n6), .C(n29), .Q(n23) );
  OAI210 U29 ( .A(n15), .B(n25), .C(n13), .Q(n30) );
  XOR30 U30 ( .A(B[11]), .B(A[11]), .C(n31), .Q(SUM[11]) );
  OAI210 U31 ( .A(n26), .B(n32), .C(n29), .Q(n31) );
  XOR20 U32 ( .A(n32), .B(n33), .Q(SUM[10]) );
  NAND20 U33 ( .A(n4), .B(n29), .Q(n33) );
  NAND20 U34 ( .A(B[10]), .B(A[10]), .Q(n29) );
  NOR20 U35 ( .A(B[10]), .B(A[10]), .Q(n26) );
  AOI210 U36 ( .A(n11), .B(n7), .C(n5), .Q(n32) );
  NAND20 U37 ( .A(B[9]), .B(A[9]), .Q(n13) );
  NOR20 U38 ( .A(B[9]), .B(A[9]), .Q(n25) );
  OAI210 U39 ( .A(n14), .B(n34), .C(n15), .Q(n11) );
  NAND20 U40 ( .A(B[8]), .B(A[8]), .Q(n15) );
  NOR20 U41 ( .A(A[8]), .B(B[8]), .Q(n34) );
  IMAJ30 U42 ( .A(B[7]), .B(n19), .C(A[7]), .Q(n14) );
  NOR20 U43 ( .A(n10), .B(n9), .Q(n19) );
endmodule


module MULT_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  input TC;
  wire   \*Logic0* , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][7] ,
         \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] ,
         \ab[6][1] , \ab[6][0] , \ab[5][7] , \ab[5][6] , \ab[5][5] ,
         \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] ,
         \ab[4][7] , \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] ,
         \ab[4][2] , \ab[4][1] , \ab[4][0] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[7][7] ,
         \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] ,
         \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][6] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][6] , \CARRYB[5][5] ,
         \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] ,
         \CARRYB[5][0] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] ,
         \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][6] ,
         \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] ,
         \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][6] , \CARRYB[1][5] ,
         \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] ,
         \CARRYB[1][0] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[7][0] ,
         \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][6] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][6] , \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] ,
         \SUMB[1][1] , ZA, ZB, \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[13] , \A2[12] , \A2[11] , \A2[10] , \A2[9] , \A2[8] ,
         \A2[7] , \A2[6] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47;
  assign ZA = A[7];
  assign ZB = B[7];

  ADD32 S14_7_0 ( .A(ZA), .B(ZB), .CI(\SUMB[7][0] ), .CO(\A2[6] ), .S(\A1[5] )
         );
  ADD32 S4_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\SUMB[7][0] ) );
  ADD32 S4_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  ADD32 S4_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  ADD32 S4_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  ADD32 S4_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  ADD32 S4_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  ADD32 S5_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\ab[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  ADD32 S14_7 ( .A(n40), .B(n32), .CI(\ab[7][7] ), .CO(\CARRYB[7][7] ), .S(
        \SUMB[7][7] ) );
  ADD32 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  ADD32 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  ADD32 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  ADD32 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  ADD32 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  ADD32 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  ADD32 S3_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\ab[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  ADD32 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  ADD32 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  ADD32 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  ADD32 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  ADD32 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  ADD32 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  ADD32 S3_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\ab[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  ADD32 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  ADD32 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  ADD32 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  ADD32 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  ADD32 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  ADD32 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  ADD32 S3_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\ab[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  ADD32 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  ADD32 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  ADD32 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  ADD32 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  ADD32 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  ADD32 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  ADD32 S3_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\ab[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  ADD32 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  ADD32 S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  ADD32 S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  ADD32 S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  ADD32 S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  ADD32 S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  ADD32 S3_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\ab[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  MULT_DW01_add_0 FS_1 ( .A({n31, \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({\A2[13] , \A2[12] , \A2[11] , \A2[10] , \A2[9] , 
        \A2[8] , \A2[7] , \A2[6] , \*Logic0* , \*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* }), .CI(\*Logic0* ), .SUM(
        PRODUCT[15:2]) );
  INV3 U2 ( .A(\ab[0][6] ), .Q(n27) );
  INV3 U3 ( .A(\ab[0][5] ), .Q(n25) );
  INV3 U4 ( .A(\ab[0][4] ), .Q(n23) );
  INV3 U5 ( .A(\ab[0][3] ), .Q(n21) );
  INV3 U6 ( .A(\ab[0][2] ), .Q(n19) );
  INV3 U7 ( .A(\ab[1][5] ), .Q(n28) );
  INV3 U8 ( .A(\ab[1][4] ), .Q(n26) );
  INV3 U9 ( .A(\ab[1][3] ), .Q(n24) );
  INV3 U10 ( .A(\ab[1][2] ), .Q(n22) );
  INV3 U11 ( .A(\ab[1][1] ), .Q(n20) );
  INV3 U12 ( .A(\ab[1][6] ), .Q(n30) );
  INV3 U13 ( .A(\CARRYB[7][7] ), .Q(n31) );
  NOR21 U14 ( .A(n15), .B(n16), .Q(\A2[13] ) );
  INV3 U15 ( .A(\ab[0][1] ), .Q(n17) );
  INV3 U16 ( .A(\ab[1][0] ), .Q(n18) );
  XOR21 U17 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Q(PRODUCT[1]) );
  INV3 U18 ( .A(\SUMB[7][7] ), .Q(n16) );
  NOR21 U19 ( .A(n27), .B(n28), .Q(\CARRYB[1][5] ) );
  XOR21 U20 ( .A(\ab[0][7] ), .B(\ab[1][6] ), .Q(\SUMB[1][6] ) );
  XOR21 U21 ( .A(\SUMB[7][1] ), .B(\CARRYB[7][0] ), .Q(\A1[6] ) );
  NOR21 U22 ( .A(n25), .B(n26), .Q(\CARRYB[1][4] ) );
  XOR21 U23 ( .A(\ab[0][6] ), .B(\ab[1][5] ), .Q(\SUMB[1][5] ) );
  NOR21 U24 ( .A(n23), .B(n24), .Q(\CARRYB[1][3] ) );
  XOR21 U25 ( .A(\ab[0][5] ), .B(\ab[1][4] ), .Q(\SUMB[1][4] ) );
  NOR21 U26 ( .A(n21), .B(n22), .Q(\CARRYB[1][2] ) );
  XOR21 U27 ( .A(\ab[0][4] ), .B(\ab[1][3] ), .Q(\SUMB[1][3] ) );
  NOR21 U28 ( .A(n19), .B(n20), .Q(\CARRYB[1][1] ) );
  XOR21 U29 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Q(\SUMB[1][2] ) );
  NOR21 U30 ( .A(n17), .B(n18), .Q(\CARRYB[1][0] ) );
  XOR21 U31 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Q(\SUMB[1][1] ) );
  INV3 U32 ( .A(\ab[0][7] ), .Q(n29) );
  XOR21 U33 ( .A(\SUMB[7][2] ), .B(\CARRYB[7][1] ), .Q(\A1[7] ) );
  NOR21 U34 ( .A(n3), .B(n4), .Q(\A2[7] ) );
  INV3 U35 ( .A(\CARRYB[7][0] ), .Q(n3) );
  INV3 U36 ( .A(\SUMB[7][1] ), .Q(n4) );
  XOR21 U37 ( .A(\SUMB[7][3] ), .B(\CARRYB[7][2] ), .Q(\A1[8] ) );
  XOR21 U38 ( .A(\SUMB[7][4] ), .B(\CARRYB[7][3] ), .Q(\A1[9] ) );
  XOR21 U39 ( .A(\SUMB[7][5] ), .B(\CARRYB[7][4] ), .Q(\A1[10] ) );
  NOR21 U40 ( .A(n5), .B(n6), .Q(\A2[8] ) );
  INV3 U41 ( .A(\CARRYB[7][1] ), .Q(n5) );
  INV3 U42 ( .A(\SUMB[7][2] ), .Q(n6) );
  NOR21 U43 ( .A(n7), .B(n8), .Q(\A2[9] ) );
  INV3 U44 ( .A(\CARRYB[7][2] ), .Q(n7) );
  INV3 U45 ( .A(\SUMB[7][3] ), .Q(n8) );
  NOR21 U46 ( .A(n9), .B(n10), .Q(\A2[10] ) );
  INV3 U47 ( .A(\CARRYB[7][3] ), .Q(n9) );
  INV3 U48 ( .A(\SUMB[7][4] ), .Q(n10) );
  XOR21 U49 ( .A(\SUMB[7][6] ), .B(\CARRYB[7][5] ), .Q(\A1[11] ) );
  NOR21 U50 ( .A(n11), .B(n12), .Q(\A2[11] ) );
  INV3 U51 ( .A(\SUMB[7][5] ), .Q(n12) );
  INV3 U52 ( .A(\CARRYB[7][4] ), .Q(n11) );
  XOR21 U53 ( .A(\SUMB[7][7] ), .B(\CARRYB[7][6] ), .Q(\A1[12] ) );
  NOR21 U54 ( .A(n13), .B(n14), .Q(\A2[12] ) );
  INV3 U55 ( .A(\SUMB[7][6] ), .Q(n14) );
  INV3 U56 ( .A(\CARRYB[7][5] ), .Q(n13) );
  INV3 U57 ( .A(\CARRYB[7][6] ), .Q(n15) );
  INV3 U58 ( .A(A[1]), .Q(n46) );
  NOR21 U59 ( .A(n29), .B(n30), .Q(\CARRYB[1][6] ) );
  INV3 U60 ( .A(B[5]), .Q(n34) );
  INV3 U61 ( .A(B[3]), .Q(n36) );
  INV3 U62 ( .A(B[6]), .Q(n33) );
  INV3 U63 ( .A(B[4]), .Q(n35) );
  INV3 U64 ( .A(A[0]), .Q(n47) );
  INV3 U65 ( .A(A[2]), .Q(n45) );
  INV3 U66 ( .A(A[3]), .Q(n44) );
  INV3 U67 ( .A(ZB), .Q(n32) );
  INV3 U68 ( .A(B[2]), .Q(n37) );
  INV3 U69 ( .A(B[0]), .Q(n39) );
  INV3 U70 ( .A(B[1]), .Q(n38) );
  INV3 U71 ( .A(A[4]), .Q(n43) );
  INV3 U72 ( .A(A[5]), .Q(n42) );
  INV3 U73 ( .A(A[6]), .Q(n41) );
  INV3 U74 ( .A(ZA), .Q(n40) );
  LOGIC0 U75 ( .Q(\*Logic0* ) );
  NOR20 U76 ( .A(n32), .B(n40), .Q(\ab[7][7] ) );
  NOR20 U77 ( .A(B[6]), .B(n40), .Q(\ab[7][6] ) );
  NOR20 U78 ( .A(B[5]), .B(n40), .Q(\ab[7][5] ) );
  NOR20 U79 ( .A(B[4]), .B(n40), .Q(\ab[7][4] ) );
  NOR20 U80 ( .A(B[3]), .B(n40), .Q(\ab[7][3] ) );
  NOR20 U81 ( .A(B[2]), .B(n40), .Q(\ab[7][2] ) );
  NOR20 U82 ( .A(B[1]), .B(n40), .Q(\ab[7][1] ) );
  NOR20 U83 ( .A(B[0]), .B(n40), .Q(\ab[7][0] ) );
  NOR20 U84 ( .A(A[6]), .B(n32), .Q(\ab[6][7] ) );
  NOR20 U85 ( .A(n41), .B(n33), .Q(\ab[6][6] ) );
  NOR20 U86 ( .A(n41), .B(n34), .Q(\ab[6][5] ) );
  NOR20 U87 ( .A(n41), .B(n35), .Q(\ab[6][4] ) );
  NOR20 U88 ( .A(n41), .B(n36), .Q(\ab[6][3] ) );
  NOR20 U89 ( .A(n41), .B(n37), .Q(\ab[6][2] ) );
  NOR20 U90 ( .A(n41), .B(n38), .Q(\ab[6][1] ) );
  NOR20 U91 ( .A(n41), .B(n39), .Q(\ab[6][0] ) );
  NOR20 U92 ( .A(A[5]), .B(n32), .Q(\ab[5][7] ) );
  NOR20 U93 ( .A(n33), .B(n42), .Q(\ab[5][6] ) );
  NOR20 U94 ( .A(n34), .B(n42), .Q(\ab[5][5] ) );
  NOR20 U95 ( .A(n35), .B(n42), .Q(\ab[5][4] ) );
  NOR20 U96 ( .A(n36), .B(n42), .Q(\ab[5][3] ) );
  NOR20 U97 ( .A(n37), .B(n42), .Q(\ab[5][2] ) );
  NOR20 U98 ( .A(n38), .B(n42), .Q(\ab[5][1] ) );
  NOR20 U99 ( .A(n39), .B(n42), .Q(\ab[5][0] ) );
  NOR20 U100 ( .A(A[4]), .B(n32), .Q(\ab[4][7] ) );
  NOR20 U101 ( .A(n33), .B(n43), .Q(\ab[4][6] ) );
  NOR20 U102 ( .A(n34), .B(n43), .Q(\ab[4][5] ) );
  NOR20 U103 ( .A(n35), .B(n43), .Q(\ab[4][4] ) );
  NOR20 U104 ( .A(n36), .B(n43), .Q(\ab[4][3] ) );
  NOR20 U105 ( .A(n37), .B(n43), .Q(\ab[4][2] ) );
  NOR20 U106 ( .A(n38), .B(n43), .Q(\ab[4][1] ) );
  NOR20 U107 ( .A(n39), .B(n43), .Q(\ab[4][0] ) );
  NOR20 U108 ( .A(A[3]), .B(n32), .Q(\ab[3][7] ) );
  NOR20 U109 ( .A(n33), .B(n44), .Q(\ab[3][6] ) );
  NOR20 U110 ( .A(n34), .B(n44), .Q(\ab[3][5] ) );
  NOR20 U111 ( .A(n35), .B(n44), .Q(\ab[3][4] ) );
  NOR20 U112 ( .A(n36), .B(n44), .Q(\ab[3][3] ) );
  NOR20 U113 ( .A(n37), .B(n44), .Q(\ab[3][2] ) );
  NOR20 U114 ( .A(n38), .B(n44), .Q(\ab[3][1] ) );
  NOR20 U115 ( .A(n39), .B(n44), .Q(\ab[3][0] ) );
  NOR20 U116 ( .A(A[2]), .B(n32), .Q(\ab[2][7] ) );
  NOR20 U117 ( .A(n33), .B(n45), .Q(\ab[2][6] ) );
  NOR20 U118 ( .A(n34), .B(n45), .Q(\ab[2][5] ) );
  NOR20 U119 ( .A(n35), .B(n45), .Q(\ab[2][4] ) );
  NOR20 U120 ( .A(n36), .B(n45), .Q(\ab[2][3] ) );
  NOR20 U121 ( .A(n37), .B(n45), .Q(\ab[2][2] ) );
  NOR20 U122 ( .A(n38), .B(n45), .Q(\ab[2][1] ) );
  NOR20 U123 ( .A(n39), .B(n45), .Q(\ab[2][0] ) );
  NOR20 U124 ( .A(A[1]), .B(n32), .Q(\ab[1][7] ) );
  NOR20 U125 ( .A(n33), .B(n46), .Q(\ab[1][6] ) );
  NOR20 U126 ( .A(n34), .B(n46), .Q(\ab[1][5] ) );
  NOR20 U127 ( .A(n35), .B(n46), .Q(\ab[1][4] ) );
  NOR20 U128 ( .A(n36), .B(n46), .Q(\ab[1][3] ) );
  NOR20 U129 ( .A(n37), .B(n46), .Q(\ab[1][2] ) );
  NOR20 U130 ( .A(n38), .B(n46), .Q(\ab[1][1] ) );
  NOR20 U131 ( .A(n39), .B(n46), .Q(\ab[1][0] ) );
  NOR20 U132 ( .A(A[0]), .B(n32), .Q(\ab[0][7] ) );
  NOR20 U133 ( .A(n33), .B(n47), .Q(\ab[0][6] ) );
  NOR20 U134 ( .A(n34), .B(n47), .Q(\ab[0][5] ) );
  NOR20 U135 ( .A(n35), .B(n47), .Q(\ab[0][4] ) );
  NOR20 U136 ( .A(n36), .B(n47), .Q(\ab[0][3] ) );
  NOR20 U137 ( .A(n37), .B(n47), .Q(\ab[0][2] ) );
  NOR20 U138 ( .A(n38), .B(n47), .Q(\ab[0][1] ) );
  NOR20 U139 ( .A(n39), .B(n47), .Q(PRODUCT[0]) );
endmodule


module MULT ( Mult_in_A, Mult_in_B, Mult_out );
  input [7:0] Mult_in_A;
  input [7:0] Mult_in_B;
  output [15:0] Mult_out;
  wire   n1;

  MULT_DW02_mult_0 mult_21 ( .A(Mult_in_B), .B(Mult_in_A), .TC(n1), .PRODUCT(
        Mult_out) );
  LOGIC1 U1 ( .Q(n1) );
endmodule


module ACCU_DW01_add_0 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [20:1] carry;

  ADD32 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADD32 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADD32 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADD32 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADD32 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADD32 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADD32 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADD32 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  INV3 U1 ( .A(n4), .Q(carry[17]) );
  NOR21 U2 ( .A(carry[16]), .B(A[16]), .Q(n4) );
  INV3 U3 ( .A(n3), .Q(carry[18]) );
  NOR21 U4 ( .A(carry[17]), .B(A[17]), .Q(n3) );
  INV3 U5 ( .A(n2), .Q(carry[19]) );
  NOR21 U6 ( .A(carry[18]), .B(A[18]), .Q(n2) );
  XOR21 U7 ( .A(n1), .B(A[20]), .Q(SUM[20]) );
  NOR21 U8 ( .A(carry[19]), .B(A[19]), .Q(n1) );
  XNR21 U9 ( .A(A[16]), .B(carry[16]), .Q(SUM[16]) );
  XNR21 U10 ( .A(A[17]), .B(carry[17]), .Q(SUM[17]) );
  XNR21 U11 ( .A(A[19]), .B(carry[19]), .Q(SUM[19]) );
  XNR21 U12 ( .A(A[18]), .B(carry[18]), .Q(SUM[18]) );
  NOR21 U13 ( .A(n5), .B(n6), .Q(carry[1]) );
  INV3 U14 ( .A(A[0]), .Q(n6) );
  INV3 U15 ( .A(B[0]), .Q(n5) );
  XOR20 U16 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
endmodule


module ACCU_DW01_add_1 ( A, B, CI, SUM, CO );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  wire   [20:1] carry;

  ADD32 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  ADD32 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADD32 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADD32 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADD32 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADD32 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADD32 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADD32 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADD32 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADD32 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADD32 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADD32 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADD32 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADD32 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADD32 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1]) );
  NOR21 U1 ( .A(n7), .B(n8), .Q(carry[17]) );
  INV3 U2 ( .A(A[16]), .Q(n8) );
  INV3 U3 ( .A(carry[16]), .Q(n7) );
  NOR21 U4 ( .A(n3), .B(n4), .Q(carry[19]) );
  INV3 U5 ( .A(A[18]), .Q(n4) );
  INV3 U6 ( .A(carry[18]), .Q(n3) );
  NOR21 U7 ( .A(n5), .B(n6), .Q(carry[18]) );
  INV3 U8 ( .A(A[17]), .Q(n6) );
  INV3 U9 ( .A(carry[17]), .Q(n5) );
  XOR21 U10 ( .A(carry[20]), .B(A[20]), .Q(SUM[20]) );
  NOR21 U11 ( .A(n1), .B(n2), .Q(carry[20]) );
  INV3 U12 ( .A(A[19]), .Q(n2) );
  INV3 U13 ( .A(carry[19]), .Q(n1) );
  XOR21 U14 ( .A(A[19]), .B(carry[19]), .Q(SUM[19]) );
  XOR21 U15 ( .A(A[18]), .B(carry[18]), .Q(SUM[18]) );
  XOR21 U16 ( .A(A[17]), .B(carry[17]), .Q(SUM[17]) );
  XOR21 U17 ( .A(A[16]), .B(carry[16]), .Q(SUM[16]) );
  XOR21 U18 ( .A(A[0]), .B(B[0]), .Q(SUM[0]) );
  NOR21 U19 ( .A(n9), .B(n10), .Q(carry[1]) );
  INV3 U20 ( .A(A[0]), .Q(n10) );
  INV3 U21 ( .A(B[0]), .Q(n9) );
endmodule


module ACCU ( CLK, RESET, Accu_in, Accu_ctrl, Accu_out );
  input [15:0] Accu_in;
  output [20:0] Accu_out;
  input CLK, RESET, Accu_ctrl;
  wire   \*Logic1* , \*Logic0* , N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n1, n2, n3, n4, n5, n6;

  DFC3 \ACCU_reg[0]  ( .D(N71), .C(CLK), .RN(n6), .Q(Accu_out[0]) );
  DFC3 \ACCU_reg[20]  ( .D(N91), .C(CLK), .RN(n6), .Q(Accu_out[20]) );
  DFC3 \ACCU_reg[1]  ( .D(N72), .C(CLK), .RN(n6), .Q(Accu_out[1]) );
  DFC3 \ACCU_reg[2]  ( .D(N73), .C(CLK), .RN(n6), .Q(Accu_out[2]) );
  DFC3 \ACCU_reg[3]  ( .D(N74), .C(CLK), .RN(n6), .Q(Accu_out[3]) );
  DFC3 \ACCU_reg[4]  ( .D(N75), .C(CLK), .RN(n6), .Q(Accu_out[4]) );
  DFC3 \ACCU_reg[5]  ( .D(N76), .C(CLK), .RN(n6), .Q(Accu_out[5]) );
  DFC3 \ACCU_reg[6]  ( .D(N77), .C(CLK), .RN(n6), .Q(Accu_out[6]) );
  DFC3 \ACCU_reg[7]  ( .D(N78), .C(CLK), .RN(n6), .Q(Accu_out[7]) );
  DFC3 \ACCU_reg[8]  ( .D(N79), .C(CLK), .RN(n6), .Q(Accu_out[8]) );
  DFC3 \ACCU_reg[9]  ( .D(N80), .C(CLK), .RN(n6), .Q(Accu_out[9]) );
  DFC3 \ACCU_reg[10]  ( .D(N81), .C(CLK), .RN(n6), .Q(Accu_out[10]) );
  DFC3 \ACCU_reg[11]  ( .D(N82), .C(CLK), .RN(n6), .Q(Accu_out[11]) );
  DFC3 \ACCU_reg[12]  ( .D(N83), .C(CLK), .RN(n6), .Q(Accu_out[12]) );
  DFC3 \ACCU_reg[13]  ( .D(N84), .C(CLK), .RN(n6), .Q(Accu_out[13]) );
  DFC3 \ACCU_reg[14]  ( .D(N85), .C(CLK), .RN(n6), .Q(Accu_out[14]) );
  DFC3 \ACCU_reg[15]  ( .D(N86), .C(CLK), .RN(n6), .Q(Accu_out[15]) );
  DFC3 \ACCU_reg[16]  ( .D(N87), .C(CLK), .RN(n6), .Q(Accu_out[16]) );
  DFC3 \ACCU_reg[17]  ( .D(N88), .C(CLK), .RN(n6), .Q(Accu_out[17]) );
  DFC3 \ACCU_reg[18]  ( .D(N89), .C(CLK), .RN(n6), .Q(Accu_out[18]) );
  DFC3 \ACCU_reg[19]  ( .D(N90), .C(CLK), .RN(n6), .Q(Accu_out[19]) );
  ACCU_DW01_add_0 add_36 ( .A(Accu_out), .B({\*Logic1* , \*Logic1* , 
        \*Logic1* , \*Logic1* , \*Logic1* , n3, Accu_in[14:0]}), .CI(
        \*Logic0* ), .SUM({N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, 
        N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29}) );
  ACCU_DW01_add_1 add_34 ( .A(Accu_out), .B({\*Logic0* , \*Logic0* , 
        \*Logic0* , \*Logic0* , \*Logic0* , n3, Accu_in[14:0]}), .CI(
        \*Logic0* ), .SUM({N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, 
        N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8}) );
  BUF2 U3 ( .A(Accu_in[15]), .Q(n3) );
  NAND22 U4 ( .A(n3), .B(n2), .Q(n8) );
  BUF2 U5 ( .A(n10), .Q(n4) );
  NOR21 U6 ( .A(n2), .B(n3), .Q(n10) );
  NOR21 U7 ( .A(n5), .B(n2), .Q(n23) );
  INV3 U8 ( .A(n3), .Q(n5) );
  INV3 U9 ( .A(n1), .Q(n2) );
  NAND31 U10 ( .A(n19), .B(n8), .C(n20), .Q(N86) );
  NAND22 U11 ( .A(N23), .B(n4), .Q(n19) );
  NAND22 U12 ( .A(N44), .B(n3), .Q(n20) );
  NAND22 U13 ( .A(n21), .B(n22), .Q(N85) );
  NAND22 U14 ( .A(Accu_in[14]), .B(n2), .Q(n22) );
  AOI221 U15 ( .A(N43), .B(n23), .C(N22), .D(n4), .Q(n21) );
  NAND22 U16 ( .A(n24), .B(n25), .Q(N84) );
  NAND22 U17 ( .A(Accu_in[13]), .B(n2), .Q(n25) );
  AOI221 U18 ( .A(N42), .B(n23), .C(N21), .D(n4), .Q(n24) );
  NAND22 U19 ( .A(n26), .B(n27), .Q(N83) );
  NAND22 U20 ( .A(Accu_in[12]), .B(n2), .Q(n27) );
  AOI221 U21 ( .A(N41), .B(n23), .C(N20), .D(n4), .Q(n26) );
  NAND22 U22 ( .A(n28), .B(n29), .Q(N82) );
  NAND22 U23 ( .A(Accu_in[11]), .B(n2), .Q(n29) );
  AOI221 U24 ( .A(N40), .B(n23), .C(N19), .D(n4), .Q(n28) );
  NAND22 U25 ( .A(n30), .B(n31), .Q(N81) );
  NAND22 U26 ( .A(Accu_in[10]), .B(n2), .Q(n31) );
  AOI221 U27 ( .A(N39), .B(n23), .C(N18), .D(n4), .Q(n30) );
  NAND22 U28 ( .A(n32), .B(n33), .Q(N80) );
  NAND22 U29 ( .A(Accu_in[9]), .B(n2), .Q(n33) );
  AOI221 U30 ( .A(N38), .B(n23), .C(N17), .D(n4), .Q(n32) );
  NAND22 U31 ( .A(n34), .B(n35), .Q(N79) );
  NAND22 U32 ( .A(Accu_in[8]), .B(n2), .Q(n35) );
  AOI221 U33 ( .A(N37), .B(n23), .C(N16), .D(n4), .Q(n34) );
  NAND22 U34 ( .A(n36), .B(n37), .Q(N78) );
  NAND22 U35 ( .A(Accu_in[7]), .B(Accu_ctrl), .Q(n37) );
  AOI221 U36 ( .A(N36), .B(n23), .C(N15), .D(n4), .Q(n36) );
  NAND22 U37 ( .A(n38), .B(n39), .Q(N77) );
  NAND22 U38 ( .A(Accu_in[6]), .B(n2), .Q(n39) );
  AOI221 U39 ( .A(N35), .B(n23), .C(N14), .D(n4), .Q(n38) );
  NAND22 U40 ( .A(n40), .B(n41), .Q(N76) );
  NAND22 U41 ( .A(Accu_in[5]), .B(n2), .Q(n41) );
  AOI221 U42 ( .A(N34), .B(n23), .C(N13), .D(n4), .Q(n40) );
  NAND22 U43 ( .A(n42), .B(n43), .Q(N75) );
  NAND22 U44 ( .A(Accu_in[4]), .B(Accu_ctrl), .Q(n43) );
  AOI221 U45 ( .A(N33), .B(n23), .C(N12), .D(n4), .Q(n42) );
  NAND22 U46 ( .A(n44), .B(n45), .Q(N74) );
  NAND22 U47 ( .A(Accu_in[3]), .B(n2), .Q(n45) );
  AOI221 U48 ( .A(N32), .B(n23), .C(N11), .D(n4), .Q(n44) );
  NAND22 U49 ( .A(n46), .B(n47), .Q(N73) );
  NAND22 U50 ( .A(Accu_in[2]), .B(n2), .Q(n47) );
  AOI221 U51 ( .A(N31), .B(n23), .C(N10), .D(n4), .Q(n46) );
  NAND22 U52 ( .A(n48), .B(n49), .Q(N72) );
  NAND22 U53 ( .A(Accu_in[1]), .B(Accu_ctrl), .Q(n49) );
  AOI221 U54 ( .A(N30), .B(n23), .C(N9), .D(n4), .Q(n48) );
  INV3 U55 ( .A(Accu_ctrl), .Q(n1) );
  NAND31 U56 ( .A(n7), .B(n8), .C(n9), .Q(N91) );
  NAND22 U57 ( .A(N28), .B(n4), .Q(n7) );
  NAND22 U58 ( .A(N49), .B(n3), .Q(n9) );
  NAND31 U59 ( .A(n11), .B(n8), .C(n12), .Q(N90) );
  NAND22 U60 ( .A(N27), .B(n4), .Q(n11) );
  NAND22 U61 ( .A(N48), .B(n3), .Q(n12) );
  NAND31 U62 ( .A(n13), .B(n8), .C(n14), .Q(N89) );
  NAND22 U63 ( .A(N26), .B(n4), .Q(n13) );
  NAND22 U64 ( .A(N47), .B(n3), .Q(n14) );
  NAND31 U65 ( .A(n15), .B(n8), .C(n16), .Q(N88) );
  NAND22 U66 ( .A(N25), .B(n4), .Q(n15) );
  NAND22 U67 ( .A(N46), .B(n3), .Q(n16) );
  NAND31 U68 ( .A(n17), .B(n8), .C(n18), .Q(N87) );
  NAND22 U69 ( .A(N24), .B(n4), .Q(n17) );
  NAND22 U70 ( .A(N45), .B(n3), .Q(n18) );
  NAND22 U71 ( .A(n50), .B(n51), .Q(N71) );
  NAND22 U72 ( .A(Accu_in[0]), .B(n2), .Q(n51) );
  AOI221 U73 ( .A(N29), .B(n23), .C(N8), .D(n4), .Q(n50) );
  INV3 U74 ( .A(RESET), .Q(n6) );
  LOGIC0 U75 ( .Q(\*Logic0* ) );
  LOGIC1 U76 ( .Q(\*Logic1* ) );
endmodule


module BUFF ( CLK, RESET, Buff_OE, Buff_in, Buff_out );
  input [7:0] Buff_in;
  output [7:0] Buff_out;
  input CLK, RESET, Buff_OE;
  wire   n1;

  DFEC1 \Buff_out_reg[7]  ( .D(Buff_in[7]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[7]) );
  DFEC1 \Buff_out_reg[6]  ( .D(Buff_in[6]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[6]) );
  DFEC1 \Buff_out_reg[5]  ( .D(Buff_in[5]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[5]) );
  DFEC1 \Buff_out_reg[4]  ( .D(Buff_in[4]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[4]) );
  DFEC1 \Buff_out_reg[3]  ( .D(Buff_in[3]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[3]) );
  DFEC1 \Buff_out_reg[2]  ( .D(Buff_in[2]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[2]) );
  DFEC1 \Buff_out_reg[1]  ( .D(Buff_in[1]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[1]) );
  DFEC1 \Buff_out_reg[0]  ( .D(Buff_in[0]), .E(Buff_OE), .C(CLK), .RN(n1), .Q(
        Buff_out[0]) );
  INV3 U2 ( .A(RESET), .Q(n1) );
endmodule


module fsm ( CLK, RESET, ADC_eoc, ADC_convst, ADC_rd, ADC_cs, DAC_wr, DAC_cs, 
        DAC_ldac, DAC_clr, Ram_Address, Delay_Line_Address, 
        Delay_Line_sample_shift, Accu_ctrl, Buff_OE );
  output [4:0] Ram_Address;
  output [4:0] Delay_Line_Address;
  input CLK, RESET, ADC_eoc;
  output ADC_convst, ADC_rd, ADC_cs, DAC_wr, DAC_cs, DAC_ldac, DAC_clr,
         Delay_Line_sample_shift, Accu_ctrl, Buff_OE;
  wire   \*Logic1* , \*Logic0* , ADC_rd, ADC_convst, N40, N43, N44, N45, N46,
         n10, n13, n15, n16, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, \add_103/carry[4] ,
         \add_103/carry[3] , \add_103/carry[2] , \Delay_Line_Address[0] , n2,
         n3, n4, n5, n6, n7, n8, n9, n11, n12, n14, n17, n38, n39;
  wire   [2:0] Current_State;
  assign DAC_clr = \*Logic1* ;
  assign DAC_ldac = \*Logic0* ;
  assign ADC_cs = ADC_rd;
  assign DAC_wr = ADC_convst;
  assign DAC_cs = ADC_convst;
  assign Delay_Line_Address[4] = Ram_Address[4];
  assign Delay_Line_Address[3] = Ram_Address[3];
  assign Delay_Line_Address[2] = Ram_Address[2];
  assign Delay_Line_Address[1] = Ram_Address[1];
  assign Delay_Line_Address[0] = \Delay_Line_Address[0] ;
  assign Ram_Address[0] = \Delay_Line_Address[0] ;

  OAI222 U3 ( .A(n15), .B(n17), .C(RESET), .D(n18), .Q(n35) );
  OAI212 U6 ( .A(RESET), .B(n5), .C(n17), .Q(n36) );
  OAI212 U7 ( .A(n15), .B(n16), .C(n21), .Q(n20) );
  OAI222 U9 ( .A(n16), .B(n17), .C(RESET), .D(n23), .Q(n37) );
  DF3 \Current_State_reg[0]  ( .D(n37), .C(CLK), .Q(Current_State[0]), .QN(n16) );
  DF3 \Current_State_reg[1]  ( .D(n35), .C(CLK), .Q(Current_State[1]), .QN(n15) );
  DF3 \Tap_Number_reg[0]  ( .D(n8), .C(CLK), .Q(\Delay_Line_Address[0] ), .QN(
        n2) );
  DF3 \Tap_Number_reg[1]  ( .D(n9), .C(CLK), .Q(Ram_Address[1]) );
  DF3 \Tap_Number_reg[2]  ( .D(n11), .C(CLK), .Q(Ram_Address[2]), .QN(n10) );
  DF3 \Tap_Number_reg[3]  ( .D(n12), .C(CLK), .Q(Ram_Address[3]) );
  DF3 \Tap_Number_reg[4]  ( .D(n14), .C(CLK), .Q(Ram_Address[4]) );
  DF3 \Current_State_reg[2]  ( .D(n36), .C(CLK), .Q(Current_State[2]), .QN(n13) );
  ADD22 \add_103/U1_1_1  ( .A(Ram_Address[1]), .B(\Delay_Line_Address[0] ), 
        .CO(\add_103/carry[2] ), .S(N43) );
  ADD22 \add_103/U1_1_2  ( .A(Ram_Address[2]), .B(\add_103/carry[2] ), .CO(
        \add_103/carry[3] ), .S(N44) );
  ADD22 \add_103/U1_1_3  ( .A(Ram_Address[3]), .B(\add_103/carry[3] ), .CO(
        \add_103/carry[4] ), .S(N45) );
  INV3 U4 ( .A(n29), .Q(n12) );
  NAND22 U5 ( .A(N45), .B(n28), .Q(n29) );
  INV3 U8 ( .A(n30), .Q(n11) );
  NAND22 U10 ( .A(N44), .B(n28), .Q(n30) );
  INV3 U11 ( .A(n31), .Q(n9) );
  NAND22 U12 ( .A(N43), .B(n28), .Q(n31) );
  INV3 U13 ( .A(n32), .Q(n8) );
  NAND22 U14 ( .A(n2), .B(n28), .Q(n32) );
  NAND22 U15 ( .A(n34), .B(n6), .Q(ADC_convst) );
  INV3 U16 ( .A(Delay_Line_sample_shift), .Q(n6) );
  NAND22 U17 ( .A(n34), .B(n24), .Q(ADC_rd) );
  NOR40 U18 ( .A(N40), .B(n10), .C(n22), .D(n33), .Q(Buff_OE) );
  NOR31 U19 ( .A(Current_State[0]), .B(Current_State[2]), .C(n15), .Q(
        Delay_Line_sample_shift) );
  NOR31 U20 ( .A(n33), .B(RESET), .C(n38), .Q(n28) );
  INV3 U21 ( .A(N40), .Q(n38) );
  INV3 U22 ( .A(n20), .Q(n5) );
  OAI311 U23 ( .A(n10), .B(N40), .C(n22), .D(Current_State[2]), .Q(n21) );
  INV3 U24 ( .A(n27), .Q(n14) );
  NAND22 U25 ( .A(N46), .B(n28), .Q(n27) );
  NAND41 U26 ( .A(Ram_Address[4]), .B(Ram_Address[3]), .C(Ram_Address[1]), .D(
        \Delay_Line_Address[0] ), .Q(n22) );
  NOR31 U27 ( .A(n16), .B(Current_State[2]), .C(n15), .Q(Accu_ctrl) );
  NOR21 U28 ( .A(Current_State[1]), .B(Current_State[0]), .Q(n26) );
  NAND22 U29 ( .A(n26), .B(Current_State[2]), .Q(n33) );
  NOR31 U30 ( .A(Current_State[1]), .B(Current_State[2]), .C(n16), .Q(n19) );
  AOI2111 U31 ( .A(ADC_eoc), .B(n19), .C(n7), .D(Delay_Line_sample_shift), .Q(
        n23) );
  INV3 U32 ( .A(n24), .Q(n7) );
  NAND22 U33 ( .A(n26), .B(n13), .Q(n24) );
  AOI211 U34 ( .A(n19), .B(n39), .C(Delay_Line_sample_shift), .Q(n18) );
  INV3 U35 ( .A(ADC_eoc), .Q(n39) );
  INV3 U36 ( .A(n25), .Q(n17) );
  NOR31 U37 ( .A(n26), .B(RESET), .C(n13), .Q(n25) );
  NOR31 U38 ( .A(n19), .B(Current_State[2]), .C(Accu_ctrl), .Q(n34) );
  LOGIC0 U39 ( .Q(\*Logic0* ) );
  LOGIC1 U40 ( .Q(\*Logic1* ) );
  XOR20 U41 ( .A(\add_103/carry[4] ), .B(Ram_Address[4]), .Q(N46) );
  NAND20 U42 ( .A(Ram_Address[4]), .B(Ram_Address[3]), .Q(n3) );
  NOR20 U43 ( .A(n2), .B(n3), .Q(n4) );
  NAND30 U44 ( .A(Ram_Address[2]), .B(Ram_Address[1]), .C(n4), .Q(N40) );
endmodule


module FILTER ( CLK, RESET, Filter_In, Filter_Out, ADC_eoc, ADC_convst, ADC_rd, 
        ADC_cs, DAC_wr, DAC_cs, DAC_ldac, DAC_clr, uC_address, uC_data_in, 
        uC_wb, uC_enable );
  input [7:0] Filter_In;
  output [7:0] Filter_Out;
  input [4:0] uC_address;
  input [7:0] uC_data_in;
  input CLK, RESET, ADC_eoc, uC_wb, uC_enable;
  output ADC_convst, ADC_rd, ADC_cs, DAC_wr, DAC_cs, DAC_ldac, DAC_clr;
  wire   Delay_Line_sample_shift, Accu_ctrl, FSM_Buff_OE, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [4:0] Delay_Line_Address;
  wire   [7:0] Delay_Line_out;
  wire   [4:0] FSM_Address;
  wire   [7:0] RAM_data_out;
  wire   [15:0] Mult_out;
  wire   [16:9] Accu_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12;

  DELAY_LINE U1 ( .RESET(RESET), .CLK(CLK), .Delay_Line_in(Filter_In), 
        .Delay_Line_address(Delay_Line_Address), .Delay_Line_sample_shift(
        Delay_Line_sample_shift), .Delay_Line_out(Delay_Line_out) );
  coeff_ram U2 ( .CLK(CLK), .RESET(RESET), .data_in(uC_data_in), .data_out(
        RAM_data_out), .address({n19, n18, n17, n16, n15}), .wb(uC_wb) );
  MULT U3 ( .Mult_in_A(Delay_Line_out), .Mult_in_B(RAM_data_out), .Mult_out(
        Mult_out) );
  ACCU U4 ( .CLK(CLK), .RESET(RESET), .Accu_in(Mult_out), .Accu_ctrl(Accu_ctrl), .Accu_out({SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, Accu_out, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12}) );
  BUFF U5 ( .CLK(CLK), .RESET(RESET), .Buff_OE(n14), .Buff_in(Accu_out), 
        .Buff_out(Filter_Out) );
  fsm U6 ( .CLK(CLK), .RESET(RESET), .ADC_eoc(ADC_eoc), .ADC_convst(ADC_convst), .ADC_rd(ADC_rd), .ADC_cs(ADC_cs), .DAC_wr(DAC_wr), .DAC_cs(DAC_cs), 
        .Ram_Address(FSM_Address), .Delay_Line_Address(Delay_Line_Address), 
        .Delay_Line_sample_shift(Delay_Line_sample_shift), .Accu_ctrl(
        Accu_ctrl), .Buff_OE(FSM_Buff_OE) );
  INV3 U21 ( .A(n12), .Q(n15) );
  AOI221 U22 ( .A(FSM_Address[0]), .B(uC_enable), .C(uC_address[0]), .D(n20), 
        .Q(n12) );
  INV3 U23 ( .A(n8), .Q(n19) );
  AOI221 U24 ( .A(uC_enable), .B(FSM_Address[4]), .C(uC_address[4]), .D(n20), 
        .Q(n8) );
  INV3 U25 ( .A(n9), .Q(n18) );
  AOI221 U26 ( .A(FSM_Address[3]), .B(uC_enable), .C(uC_address[3]), .D(n20), 
        .Q(n9) );
  INV3 U27 ( .A(n10), .Q(n17) );
  AOI221 U28 ( .A(FSM_Address[2]), .B(uC_enable), .C(uC_address[2]), .D(n20), 
        .Q(n10) );
  INV3 U29 ( .A(n11), .Q(n16) );
  AOI221 U30 ( .A(FSM_Address[1]), .B(uC_enable), .C(uC_address[1]), .D(n20), 
        .Q(n11) );
  INV3 U31 ( .A(n13), .Q(n14) );
  NAND22 U32 ( .A(FSM_Buff_OE), .B(uC_enable), .Q(n13) );
  INV3 U33 ( .A(uC_enable), .Q(n20) );
  LOGIC1 U34 ( .Q(DAC_clr) );
  LOGIC0 U35 ( .Q(DAC_ldac) );
endmodule

